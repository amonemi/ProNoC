#name:2SNs-RND1
11.5275194222563 56
10.4719324391456 52
8.83542552968544 43
7.42298150852438 37
5.51083348579494 32
4.39188837673891 31
3.63869899916381 30
2.70002048865441 28
2.14096142818721 28
1.51590314324332 27
1.17545096574806 27
0.807304769028575 27


#name:4SNs-RND1
11.7943266379455 53
10.7802507035047 48
8.99547665784757 40
7.521492526665  34
5.56633023286496 29
4.40880089387342 28
3.64222985213686 28
2.70002048865441 27
2.14096142818721 27
1.51590314324332 27
1.17545096574806 27
0.807304769028575 27

