#name:XY
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:WEST_FIRST
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:NORTH_LAST
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:NEGETIVE_FIRST
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:DUATO_NORTH_LAST1$
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:DUATO_NORTH_LAST2$
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:DUATO_NORTH_LAST3$
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:DUATO_XY1$
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:DUATO_XY2$
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:DUATO_XY3$
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:XY
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:WEST_FIRST
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:NORTH_LAST
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:NEGETIVE_FIRST
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:DUATO_NORTH_LAST1$
47.980455 38.708594


#name:DUATO_NORTH_LAST2$
47.980455 38.708594


#name:DUATO_NORTH_LAST3$
47.980455 38.708594


#name:DUATO_XY1$
47.980455 38.708594


#name:DUATO_XY2$
47.980455 38.708594


#name:DUATO_XY3$
47.980455 38.708594


#name:XY
#name:XY
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:WEST_FIRST
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:NORTH_LAST
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:NEGETIVE_FIRST
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:DUATO_NORTH_LAST1$
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:DUATO_NORTH_LAST2$
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:DUATO_NORTH_LAST3$
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:DUATO_XY1$
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:DUATO_XY2$
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:DUATO_XY3$
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:XY
32.287126 35.967969
29.429231 33.947656
25.710582 32.522656
27.103751 25.796094
25.289253 19.316406
20.643614 14.332031
17.258680 14.875781
12.996676 14.790625
10.422825 12.989844
5.815840 14.262500


#name:WEST_FIRST
32.287126 35.967969
29.429231 33.947656
25.710582 32.522656
27.103751 25.796094
25.289253 19.316406
20.643614 14.332031
17.258680 14.875781
12.996676 14.790625
10.422825 12.989844
5.815840 14.262500


#name:NORTH_LAST
32.287126 35.967969
29.429231 33.947656
25.710582 32.522656
27.103751 25.796094
25.289253 19.316406
20.643614 14.332031
17.258680 14.875781
12.996676 14.790625
10.422825 12.989844
5.815840 14.262500


#name:NEGETIVE_FIRST
32.287126 35.967969
29.429231 33.947656
25.710582 32.522656
27.103751 25.796094
25.289253 19.316406
20.643614 14.332031
17.258680 14.875781
12.996676 14.790625
10.422825 12.989844
5.815840 14.262500


#name:DUATO_NORTH_LAST1$
32.287126 35.967969
29.429231 33.947656
25.710582 32.522656
27.103751 25.796094
25.289253 19.316406
20.643614 14.332031
17.258680 14.875781
12.996676 14.790625
10.422825 12.989844
5.815840 14.262500


#name:DUATO_NORTH_LAST2$
32.287126 35.967969
29.429231 33.947656
25.710582 32.522656
27.103751 25.796094
25.289253 19.316406
20.643614 14.332031
17.258680 14.875781
12.996676 14.790625
10.422825 12.989844
5.815840 14.262500


#name:DUATO_NORTH_LAST3$
32.287126 35.967969
29.429231 33.947656
25.710582 32.522656
27.103751 25.796094
25.289253 19.316406
20.643614 14.332031
17.258680 14.875781
12.996676 14.790625
10.422825 12.989844
5.815840 14.262500


#name:DUATO_XY1$
32.287126 35.967969
29.429231 33.947656
25.710582 32.522656
27.103751 25.796094
25.289253 19.316406
20.643614 14.332031
17.258680 14.875781
12.996676 14.790625
10.422825 12.989844
5.815840 14.262500


#name:DUATO_XY2$
32.287126 35.967969
29.429231 33.947656
25.710582 32.522656
27.103751 25.796094
25.289253 19.316406
20.643614 14.332031
17.258680 14.875781
12.996676 14.790625
10.422825 12.989844
5.815840 14.262500


#name:DUATO_XY3$
32.287126 35.967969
29.429231 33.947656
25.710582 32.522656
27.103751 25.796094
25.289253 19.316406
20.643614 14.332031
17.258680 14.875781
12.996676 14.790625
10.422825 12.989844
5.815840 14.262500


