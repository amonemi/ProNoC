36.311782 75.779156
36.220264 70.454937
33.946492 67.630938
34.101081 60.286844
35.151573 43.044219
29.917540 16.072063
24.951008 14.320156
18.731780 13.402656
14.994330 13.330312
8.338994 13.229281


36.022649 77.251563
35.165350 71.876094
34.507549 68.080906
34.026867 60.488375
34.884862 43.689250
29.917540 16.099250
24.951008 14.329281
18.731780 13.390219
14.994330 13.315781
8.338994 13.217500
