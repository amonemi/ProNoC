#name:XY
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:WEST_FIRST
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:NORTH_LAST
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438


#name:NEGETIVE_FIRST
47.980455 38.708594
40.151965 25.397656
33.659488 20.351562
29.249006 15.997656
25.680525 14.021094
20.643614 13.086719
17.258680 13.425000
12.996676 13.765625
10.422825 12.707812
5.815840 13.698438
