module JTAGB (
         output JTCK,
         output JRTI1,
         output JRTI2,
         output JTDI,
         output JSHIFT,
         output JUPDATE,
         output JRSTN,
         output JCE1,
         output JCE2,
         input JTDO1,
         input JTDO2
      ) /*synthesis syn_black_box */; 
      
endmodule
