`include "system_conf.v"

`timescale 1 ns / 1 ps
module lm32_monitor_ram (DataInA, DataInB, AddressA, AddressB, ClockA, 
			 ClockB, ClockEnA, ClockEnB, WrA, WrB, ResetA, ResetB, QA, QB);
   input [31:0] DataInA;
   input [31:0] DataInB;
   input [8:0] 	AddressA;
   input [8:0] 	AddressB;
   input 	ClockA;
   input 	ClockB;
   input 	ClockEnA;
   input 	ClockEnB;
   input 	WrA;
   input 	WrB;
   input 	ResetA;
   input 	ResetB;
   output [31:0] QA;
   output [31:0] QB;

   parameter 	 lat_family = `LATTICE_FAMILY;
   
   generate
      if (lat_family == "EC" || lat_family == "ECP" || lat_family == "XP") begin
	 /* Verilog netlist generated by SCUBA ispLever_v51_SP2_Build (10) */
	 /* Module Version: 2.0 */
	 /* c:\applications\ispTools5.1\ispfpga\bin\nt\scuba.exe -w -lang verilog -synth synplify -bus_exp 7 -bb -arch ep5g00 -type bram -wp 11 -rp 1010 -addr_width 9 -data_width 32 -num_rows 512 -gsr ENABLED -writemode NORMAL -resetmode ASYNC -memfile ../../source/jtag_rom_monitor/rom.mem -memformat hex  */
	 
	 // synopsys translate_off
	 defparam lm32_monitor_ram_0_0_1.INITVAL_1F = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_1E = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_1D = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_1C = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_1B = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_1A = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_19 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_18 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_17 = 320'h00000000000000000000000000000000000000003FF8C300003FF8E300003FF90300003FF923FF5B;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_16 = 320'h1004F3FF95300003FF97300003FF99300003FF9B300003FF9D300003FF9F300003FFA1300003FFFB;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_15 = 320'h0000130001100003FF691001400000068003FF7E058003FF803FFFB300013FF7800001100001FFB3;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_14 = 320'h00000068003FF89058003FF8B3FFB93FF9B008003FFBC300000FFBE1001B000331001A0002C10019;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_13 = 320'h00035100180003510013000301001200030100110003010010000301000900030100080003010007;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_12 = 320'h010003FF97058003FFAA3FFFC00800078003FFDB3FFBD0080000004100063FFA2000000001C10004;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_11 = 320'h000083000C2001010014000183001C0000000000000001000000000000000000010000100010FFF3;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_10 = 320'h10063000481004D0003F1006D0003E1007200024100570001D10077010003FFC210000100540FFFF;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_0F = 320'h0080010000100540FFFF008000700010004000083000C2001010014000183001C0FFE40000000008;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_0E = 320'h100043FFDD100083FFDF100093FFE11000A3FFE31000B10008100040FFF8000000000C1000410008;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_0D = 320'h100083FFE7100093FFE91000A3FFEB1000B3FFED100040FFF400000200000FFFF010000000000002;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_0C = 320'h10054100000FFFF01000100FF00000100FF000000FFFE10100010000000000070300803000030090;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_0B = 320'h300003008C300003008820078100743006C2006810064000603005C2005810054000503004C20048;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_0A = 320'h10044000403003C2003810034000303002C2002810024000203001C2001810014000103000C20008;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_09 = 320'h100040000000070200802000020090200002008C20000200883007C100743006C200681006400060;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_08 = 320'h3005C2005810054000503004C2004810044000403003C2003810034000303002C200281002400020;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_07 = 320'h3001C2001810014000103000C2000810004000001F9940E000000001007410000100841000110001;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_06 = 320'h100011000110001100FF1F99410090008001008C0080010088008003007C20078000703006C20068;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_05 = 320'h10064000603005C2005810054000503004C2004810044000403003C2003810034000303002C20028;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_04 = 320'h10024000203001C2001810014000103000C200081000400000000001066C3FFC530000007F40E000;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_03 = 320'h000000003B000B500800200800000A00000000000000000043000BD0080020080000120000000000;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_02 = 320'h000000004B000C500800200800001A00000000000000000053000CD0080020080000220000000000;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_01 = 320'h0000000081000D500800300800002A00000000000000000063000DD0080020080000320000000000;
	 defparam lm32_monitor_ram_0_0_1.INITVAL_00 = 320'h0000000091000E500800300800003A00000000000000000000000000000000000000000003F00000;
	 defparam lm32_monitor_ram_0_0_1.CSDECODE_B = "000";
	 defparam lm32_monitor_ram_0_0_1.CSDECODE_A = "000";
	 defparam lm32_monitor_ram_0_0_1.WRITEMODE_B = "NORMAL";
	 defparam lm32_monitor_ram_0_0_1.WRITEMODE_A = "NORMAL";
	 defparam lm32_monitor_ram_0_0_1.GSR = "ENABLED";
	 defparam lm32_monitor_ram_0_0_1.RESETMODE = "ASYNC";
	 defparam lm32_monitor_ram_0_0_1.REGMODE_B = "NOREG";
	 defparam lm32_monitor_ram_0_0_1.REGMODE_A = "NOREG";
	 defparam lm32_monitor_ram_0_0_1.DATA_WIDTH_B = 18;
	 defparam lm32_monitor_ram_0_0_1.DATA_WIDTH_A = 18;
	 // synopsys translate_on
	 DP8KA lm32_monitor_ram_0_0_1 (.CEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), 
				       .CSA0(scuba_vlo), .CSA1(scuba_vlo), .CSA2(scuba_vlo), .RSTA(ResetA), 
				       .CEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB0(scuba_vlo), .CSB1(scuba_vlo), 
				       .CSB2(scuba_vlo), .RSTB(ResetB), .DIA0(DataInA[0]), .DIA1(DataInA[1]), 
				       .DIA2(DataInA[2]), .DIA3(DataInA[3]), .DIA4(DataInA[4]), .DIA5(DataInA[5]), 
				       .DIA6(DataInA[6]), .DIA7(DataInA[7]), .DIA8(DataInA[8]), .DIA9(DataInA[9]), 
				       .DIA10(DataInA[10]), .DIA11(DataInA[11]), .DIA12(DataInA[12]), .DIA13(DataInA[13]), 
				       .DIA14(DataInA[14]), .DIA15(DataInA[15]), .DIA16(DataInA[16]), .DIA17(DataInA[17]), 
				       .ADA0(scuba_vhi), .ADA1(scuba_vhi), .ADA2(scuba_vlo), .ADA3(scuba_vlo), 
				       .ADA4(AddressA[0]), .ADA5(AddressA[1]), .ADA6(AddressA[2]), .ADA7(AddressA[3]), 
				       .ADA8(AddressA[4]), .ADA9(AddressA[5]), .ADA10(AddressA[6]), .ADA11(AddressA[7]), 
				       .ADA12(AddressA[8]), .DIB0(DataInB[0]), .DIB1(DataInB[1]), .DIB2(DataInB[2]), 
				       .DIB3(DataInB[3]), .DIB4(DataInB[4]), .DIB5(DataInB[5]), .DIB6(DataInB[6]), 
				       .DIB7(DataInB[7]), .DIB8(DataInB[8]), .DIB9(DataInB[9]), .DIB10(DataInB[10]), 
				       .DIB11(DataInB[11]), .DIB12(DataInB[12]), .DIB13(DataInB[13]), .DIB14(DataInB[14]), 
				       .DIB15(DataInB[15]), .DIB16(DataInB[16]), .DIB17(DataInB[17]), .ADB0(scuba_vhi), 
				       .ADB1(scuba_vhi), .ADB2(scuba_vlo), .ADB3(scuba_vlo), .ADB4(AddressB[0]), 
				       .ADB5(AddressB[1]), .ADB6(AddressB[2]), .ADB7(AddressB[3]), .ADB8(AddressB[4]), 
				       .ADB9(AddressB[5]), .ADB10(AddressB[6]), .ADB11(AddressB[7]), .ADB12(AddressB[8]), 
				       .DOA0(QA[0]), .DOA1(QA[1]), .DOA2(QA[2]), .DOA3(QA[3]), .DOA4(QA[4]), 
				       .DOA5(QA[5]), .DOA6(QA[6]), .DOA7(QA[7]), .DOA8(QA[8]), .DOA9(QA[9]), 
				       .DOA10(QA[10]), .DOA11(QA[11]), .DOA12(QA[12]), .DOA13(QA[13]), 
				       .DOA14(QA[14]), .DOA15(QA[15]), .DOA16(QA[16]), .DOA17(QA[17]), 
				       .DOB0(QB[0]), .DOB1(QB[1]), .DOB2(QB[2]), .DOB3(QB[3]), .DOB4(QB[4]), 
				       .DOB5(QB[5]), .DOB6(QB[6]), .DOB7(QB[7]), .DOB8(QB[8]), .DOB9(QB[9]), 
				       .DOB10(QB[10]), .DOB11(QB[11]), .DOB12(QB[12]), .DOB13(QB[13]), 
				       .DOB14(QB[14]), .DOB15(QB[15]), .DOB16(QB[16]), .DOB17(QB[17]))
           /* synthesis INITVAL_1F="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1E="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1D="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1C="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1B="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1A="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_19="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_18="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_17="0x00000000000000000000000000000000000000003FF8C300003FF8E300003FF90300003FF923FF5B" */
           /* synthesis INITVAL_16="0x1004F3FF95300003FF97300003FF99300003FF9B300003FF9D300003FF9F300003FFA1300003FFFB" */
           /* synthesis INITVAL_15="0x0000130001100003FF691001400000068003FF7E058003FF803FFFB300013FF7800001100001FFB3" */
           /* synthesis INITVAL_14="0x00000068003FF89058003FF8B3FFB93FF9B008003FFBC300000FFBE1001B000331001A0002C10019" */
           /* synthesis INITVAL_13="0x00035100180003510013000301001200030100110003010010000301000900030100080003010007" */
           /* synthesis INITVAL_12="0x010003FF97058003FFAA3FFFC00800078003FFDB3FFBD0080000004100063FFA2000000001C10004" */
           /* synthesis INITVAL_11="0x000083000C2001010014000183001C0000000000000001000000000000000000010000100010FFF3" */
           /* synthesis INITVAL_10="0x10063000481004D0003F1006D0003E1007200024100570001D10077010003FFC210000100540FFFF" */
           /* synthesis INITVAL_0F="0x0080010000100540FFFF008000700010004000083000C2001010014000183001C0FFE40000000008" */
           /* synthesis INITVAL_0E="0x100043FFDD100083FFDF100093FFE11000A3FFE31000B10008100040FFF8000000000C1000410008" */
           /* synthesis INITVAL_0D="0x100083FFE7100093FFE91000A3FFEB1000B3FFED100040FFF400000200000FFFF010000000000002" */
           /* synthesis INITVAL_0C="0x10054100000FFFF01000100FF00000100FF000000FFFE10100010000000000070300803000030090" */
           /* synthesis INITVAL_0B="0x300003008C300003008820078100743006C2006810064000603005C2005810054000503004C20048" */
           /* synthesis INITVAL_0A="0x10044000403003C2003810034000303002C2002810024000203001C2001810014000103000C20008" */
           /* synthesis INITVAL_09="0x100040000000070200802000020090200002008C20000200883007C100743006C200681006400060" */
           /* synthesis INITVAL_08="0x3005C2005810054000503004C2004810044000403003C2003810034000303002C200281002400020" */
           /* synthesis INITVAL_07="0x3001C2001810014000103000C2000810004000001F9940E000000001007410000100841000110001" */
           /* synthesis INITVAL_06="0x100011000110001100FF1F99410090008001008C0080010088008003007C20078000703006C20068" */
           /* synthesis INITVAL_05="0x10064000603005C2005810054000503004C2004810044000403003C2003810034000303002C20028" */
           /* synthesis INITVAL_04="0x10024000203001C2001810014000103000C200081000400000000001066C3FFC530000007F40E000" */
           /* synthesis INITVAL_03="0x000000003B000B500800200800000A00000000000000000043000BD0080020080000120000000000" */
           /* synthesis INITVAL_02="0x000000004B000C500800200800001A00000000000000000053000CD0080020080000220000000000" */
           /* synthesis INITVAL_01="0x0000000081000D500800300800002A00000000000000000063000DD0080020080000320000000000" */
           /* synthesis INITVAL_00="0x0000000091000E500800300800003A00000000000000000000000000000000000000000003F00000" */
           /* synthesis CSDECODE_B="000" */
           /* synthesis CSDECODE_A="000" */
           /* synthesis WRITEMODE_B="NORMAL" */
           /* synthesis WRITEMODE_A="NORMAL" */
           /* synthesis GSR="ENABLED" */
           /* synthesis RESETMODE="ASYNC" */
           /* synthesis REGMODE_B="NOREG" */
           /* synthesis REGMODE_A="NOREG" */
           /* synthesis DATA_WIDTH_B="18" */
           /* synthesis DATA_WIDTH_A="18" */;

	 VHI scuba_vhi_inst (.Z(scuba_vhi));

	 VLO scuba_vlo_inst (.Z(scuba_vlo));

	 // synopsys translate_off
	 defparam lm32_monitor_ram_0_1_0.INITVAL_1F = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_1E = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_1D = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_1C = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_1B = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_1A = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_19 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_18 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_17 = 320'h0000000000000000000000000000000000000000038FF034D2038FF034C2038FF0349A038FF03EFF;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_16 = 320'h00D00038FF034CA038FF03492038FF0348A038FF03482038FF0344A038FF03442038FF0343A038FF;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_15 = 320'h00D6300D5A00C5803EFF0136300D0302E0803EFF02E0803EFF038FF00D5A03EFF00D630105801363;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_14 = 320'h00D0302E0803EFF02E0803EFF038FF03EFF02E70038FF034DA0170801F100110801F100110801F10;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_13 = 320'h0110801F100110801F100110801F100110801F100110801F100110801F100110801F100110801F08;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_12 = 320'h02E0803EFF02E0803EFF038FF02E7802430038FF03EFF02E780110801F0803EFF030E800DE700AE7;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_11 = 320'h00AE400AE300AE300AE300AE300AE200D0000D0000D000342000D0000D0000D000341800D0001708;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_10 = 320'h01F100110801F100110801F100110801F100110801F100110801F0802E0803EFF0347000D0001708;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_0F = 320'h024700347000D00017080247002E08016E7016E4016E3016E3016E3016E3016E200DE7030E800DE7;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_0E = 320'h00AE703EFF010E003EFF010E003EFF010E003EFF010E0016E0016E700DE7030E800DE700AE700AE0;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_0D = 320'h00CE003EFF00CE003EFF00CE003EFF00CE003EFF016E700DE7030E8034700171002470030E801108;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_0C = 320'h01F0803470017100247000808030E80081003478011080081002478030F800AE700AE70340700AE7;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_0B = 320'h0344F00AE70343F00AE700AE700AE700AE600AE600AE600AE600AE500AE500AE500AE500AE400AE4;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_0A = 320'h00AE400AE400AE300AE300AE300AE300AE200AE200AE200AE200AE100AE100AE100AE100AE000AE0;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_09 = 320'h00AE0030F000AE700AE70340700AE70344F00AE70343F00AE700AE700AE700AE600AE600AE600AE6;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_08 = 320'h00AE500AE500AE500AE500AE400AE400AE400AE400AE300AE300AE300AE300AE200AE200AE200AE2;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_07 = 320'h00AE100AE100AE100AE100AE000AE000AE0030E800DEF02EE8016E8016E800AE8016E80000800008;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_06 = 320'h0000800008000080080800DE8016E802400016E802448016E802438016EF016EF016EF016EE016EE;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_05 = 320'h016EE016EE016ED016ED016ED016ED016EC016EC016EC016EC016EB016EB016EB016EB016EA016EA;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_04 = 320'h016EA016EA016E9016E9016E9016E9016E8016E8016E802600016E800DEF038FF00D0700DE702EE8;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_03 = 320'h00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_02 = 320'h00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_01 = 320'h00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600;
	 defparam lm32_monitor_ram_0_1_0.INITVAL_00 = 320'h00D000380003E0002EE0016E703E0002EE80260000D0000D0000D0000D0000D0000D0003E0002600;
	 defparam lm32_monitor_ram_0_1_0.CSDECODE_B = "000";
	 defparam lm32_monitor_ram_0_1_0.CSDECODE_A = "000";
	 defparam lm32_monitor_ram_0_1_0.WRITEMODE_B = "NORMAL";
	 defparam lm32_monitor_ram_0_1_0.WRITEMODE_A = "NORMAL";
	 defparam lm32_monitor_ram_0_1_0.GSR = "ENABLED";
	 defparam lm32_monitor_ram_0_1_0.RESETMODE = "ASYNC";
	 defparam lm32_monitor_ram_0_1_0.REGMODE_B = "NOREG";
	 defparam lm32_monitor_ram_0_1_0.REGMODE_A = "NOREG";
	 defparam lm32_monitor_ram_0_1_0.DATA_WIDTH_B = 18;
	 defparam lm32_monitor_ram_0_1_0.DATA_WIDTH_A = 18;
	 // synopsys translate_on
	 DP8KA lm32_monitor_ram_0_1_0 (.CEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), 
				       .CSA0(scuba_vlo), .CSA1(scuba_vlo), .CSA2(scuba_vlo), .RSTA(ResetA), 
				       .CEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB0(scuba_vlo), .CSB1(scuba_vlo), 
				       .CSB2(scuba_vlo), .RSTB(ResetB), .DIA0(DataInA[18]), .DIA1(DataInA[19]), 
				       .DIA2(DataInA[20]), .DIA3(DataInA[21]), .DIA4(DataInA[22]), .DIA5(DataInA[23]), 
				       .DIA6(DataInA[24]), .DIA7(DataInA[25]), .DIA8(DataInA[26]), .DIA9(DataInA[27]), 
				       .DIA10(DataInA[28]), .DIA11(DataInA[29]), .DIA12(DataInA[30]), .DIA13(DataInA[31]), 
				       .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), .DIA17(scuba_vlo), 
				       .ADA0(scuba_vhi), .ADA1(scuba_vhi), .ADA2(scuba_vlo), .ADA3(scuba_vlo), 
				       .ADA4(AddressA[0]), .ADA5(AddressA[1]), .ADA6(AddressA[2]), .ADA7(AddressA[3]), 
				       .ADA8(AddressA[4]), .ADA9(AddressA[5]), .ADA10(AddressA[6]), .ADA11(AddressA[7]), 
				       .ADA12(AddressA[8]), .DIB0(DataInB[18]), .DIB1(DataInB[19]), .DIB2(DataInB[20]), 
				       .DIB3(DataInB[21]), .DIB4(DataInB[22]), .DIB5(DataInB[23]), .DIB6(DataInB[24]), 
				       .DIB7(DataInB[25]), .DIB8(DataInB[26]), .DIB9(DataInB[27]), .DIB10(DataInB[28]), 
				       .DIB11(DataInB[29]), .DIB12(DataInB[30]), .DIB13(DataInB[31]), .DIB14(scuba_vlo), 
				       .DIB15(scuba_vlo), .DIB16(scuba_vlo), .DIB17(scuba_vlo), .ADB0(scuba_vhi), 
				       .ADB1(scuba_vhi), .ADB2(scuba_vlo), .ADB3(scuba_vlo), .ADB4(AddressB[0]), 
				       .ADB5(AddressB[1]), .ADB6(AddressB[2]), .ADB7(AddressB[3]), .ADB8(AddressB[4]), 
				       .ADB9(AddressB[5]), .ADB10(AddressB[6]), .ADB11(AddressB[7]), .ADB12(AddressB[8]), 
				       .DOA0(QA[18]), .DOA1(QA[19]), .DOA2(QA[20]), .DOA3(QA[21]), .DOA4(QA[22]), 
				       .DOA5(QA[23]), .DOA6(QA[24]), .DOA7(QA[25]), .DOA8(QA[26]), .DOA9(QA[27]), 
				       .DOA10(QA[28]), .DOA11(QA[29]), .DOA12(QA[30]), .DOA13(QA[31]), 
				       .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(QB[18]), .DOB1(QB[19]), 
				       .DOB2(QB[20]), .DOB3(QB[21]), .DOB4(QB[22]), .DOB5(QB[23]), .DOB6(QB[24]), 
				       .DOB7(QB[25]), .DOB8(QB[26]), .DOB9(QB[27]), .DOB10(QB[28]), .DOB11(QB[29]), 
				       .DOB12(QB[30]), .DOB13(QB[31]), .DOB14(), .DOB15(), .DOB16(), .DOB17())
           /* synthesis INITVAL_1F="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1E="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1D="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1C="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1B="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1A="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_19="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_18="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_17="0x0000000000000000000000000000000000000000038FF034D2038FF034C2038FF0349A038FF03EFF" */
           /* synthesis INITVAL_16="0x00D00038FF034CA038FF03492038FF0348A038FF03482038FF0344A038FF03442038FF0343A038FF" */
           /* synthesis INITVAL_15="0x00D6300D5A00C5803EFF0136300D0302E0803EFF02E0803EFF038FF00D5A03EFF00D630105801363" */
           /* synthesis INITVAL_14="0x00D0302E0803EFF02E0803EFF038FF03EFF02E70038FF034DA0170801F100110801F100110801F10" */
           /* synthesis INITVAL_13="0x0110801F100110801F100110801F100110801F100110801F100110801F100110801F100110801F08" */
           /* synthesis INITVAL_12="0x02E0803EFF02E0803EFF038FF02E7802430038FF03EFF02E780110801F0803EFF030E800DE700AE7" */
           /* synthesis INITVAL_11="0x00AE400AE300AE300AE300AE300AE200D0000D0000D000342000D0000D0000D000341800D0001708" */
           /* synthesis INITVAL_10="0x01F100110801F100110801F100110801F100110801F100110801F0802E0803EFF0347000D0001708" */
           /* synthesis INITVAL_0F="0x024700347000D00017080247002E08016E7016E4016E3016E3016E3016E3016E200DE7030E800DE7" */
           /* synthesis INITVAL_0E="0x00AE703EFF010E003EFF010E003EFF010E003EFF010E0016E0016E700DE7030E800DE700AE700AE0" */
           /* synthesis INITVAL_0D="0x00CE003EFF00CE003EFF00CE003EFF00CE003EFF016E700DE7030E8034700171002470030E801108" */
           /* synthesis INITVAL_0C="0x01F0803470017100247000808030E80081003478011080081002478030F800AE700AE70340700AE7" */
           /* synthesis INITVAL_0B="0x0344F00AE70343F00AE700AE700AE700AE600AE600AE600AE600AE500AE500AE500AE500AE400AE4" */
           /* synthesis INITVAL_0A="0x00AE400AE400AE300AE300AE300AE300AE200AE200AE200AE200AE100AE100AE100AE100AE000AE0" */
           /* synthesis INITVAL_09="0x00AE0030F000AE700AE70340700AE70344F00AE70343F00AE700AE700AE700AE600AE600AE600AE6" */
           /* synthesis INITVAL_08="0x00AE500AE500AE500AE500AE400AE400AE400AE400AE300AE300AE300AE300AE200AE200AE200AE2" */
           /* synthesis INITVAL_07="0x00AE100AE100AE100AE100AE000AE000AE0030E800DEF02EE8016E8016E800AE8016E80000800008" */
           /* synthesis INITVAL_06="0x0000800008000080080800DE8016E802400016E802448016E802438016EF016EF016EF016EE016EE" */
           /* synthesis INITVAL_05="0x016EE016EE016ED016ED016ED016ED016EC016EC016EC016EC016EB016EB016EB016EB016EA016EA" */
           /* synthesis INITVAL_04="0x016EA016EA016E9016E9016E9016E9016E8016E8016E802600016E800DEF038FF00D0700DE702EE8" */
           /* synthesis INITVAL_03="0x00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600" */
           /* synthesis INITVAL_02="0x00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600" */
           /* synthesis INITVAL_01="0x00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600" */
           /* synthesis INITVAL_00="0x00D000380003E0002EE0016E703E0002EE80260000D0000D0000D0000D0000D0000D0003E0002600" */
           /* synthesis CSDECODE_B="000" */
           /* synthesis CSDECODE_A="000" */
           /* synthesis WRITEMODE_B="NORMAL" */
           /* synthesis WRITEMODE_A="NORMAL" */
           /* synthesis GSR="ENABLED" */
           /* synthesis RESETMODE="ASYNC" */
           /* synthesis REGMODE_B="NOREG" */
           /* synthesis REGMODE_A="NOREG" */
           /* synthesis DATA_WIDTH_B="18" */
           /* synthesis DATA_WIDTH_A="18" */;



	 // exemplar begin
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_1F 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_1E 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_1D 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_1C 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_1B 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_1A 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_19 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_18 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_17 0x00000000000000000000000000000000000000003FF8C300003FF8E300003FF90300003FF923FF5B
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_16 0x1004F3FF95300003FF97300003FF99300003FF9B300003FF9D300003FF9F300003FFA1300003FFFB
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_15 0x0000130001100003FF691001400000068003FF7E058003FF803FFFB300013FF7800001100001FFB3
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_14 0x00000068003FF89058003FF8B3FFB93FF9B008003FFBC300000FFBE1001B000331001A0002C10019
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_13 0x00035100180003510013000301001200030100110003010010000301000900030100080003010007
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_12 0x010003FF97058003FFAA3FFFC00800078003FFDB3FFBD0080000004100063FFA2000000001C10004
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_11 0x000083000C2001010014000183001C0000000000000001000000000000000000010000100010FFF3
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_10 0x10063000481004D0003F1006D0003E1007200024100570001D10077010003FFC210000100540FFFF
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_0F 0x0080010000100540FFFF008000700010004000083000C2001010014000183001C0FFE40000000008
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_0E 0x100043FFDD100083FFDF100093FFE11000A3FFE31000B10008100040FFF8000000000C1000410008
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_0D 0x100083FFE7100093FFE91000A3FFEB1000B3FFED100040FFF400000200000FFFF010000000000002
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_0C 0x10054100000FFFF01000100FF00000100FF000000FFFE10100010000000000070300803000030090
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_0B 0x300003008C300003008820078100743006C2006810064000603005C2005810054000503004C20048
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_0A 0x10044000403003C2003810034000303002C2002810024000203001C2001810014000103000C20008
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_09 0x100040000000070200802000020090200002008C20000200883007C100743006C200681006400060
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_08 0x3005C2005810054000503004C2004810044000403003C2003810034000303002C200281002400020
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_07 0x3001C2001810014000103000C2000810004000001F9940E000000001007410000100841000110001
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_06 0x100011000110001100FF1F99410090008001008C0080010088008003007C20078000703006C20068
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_05 0x10064000603005C2005810054000503004C2004810044000403003C2003810034000303002C20028
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_04 0x10024000203001C2001810014000103000C200081000400000000001066C3FFC530000007F40E000
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_03 0x000000003B000B500800200800000A00000000000000000043000BD0080020080000120000000000
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_02 0x000000004B000C500800200800001A00000000000000000053000CD0080020080000220000000000
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_01 0x0000000081000D500800300800002A00000000000000000063000DD0080020080000320000000000
	 // exemplar attribute lm32_monitor_ram_0_0_1 INITVAL_00 0x0000000091000E500800300800003A00000000000000000000000000000000000000000003F00000
	 // exemplar attribute lm32_monitor_ram_0_0_1 CSDECODE_B 000
	 // exemplar attribute lm32_monitor_ram_0_0_1 CSDECODE_A 000
	 // exemplar attribute lm32_monitor_ram_0_0_1 WRITEMODE_B NORMAL
	 // exemplar attribute lm32_monitor_ram_0_0_1 WRITEMODE_A NORMAL
	 // exemplar attribute lm32_monitor_ram_0_0_1 GSR ENABLED
	 // exemplar attribute lm32_monitor_ram_0_0_1 RESETMODE ASYNC
	 // exemplar attribute lm32_monitor_ram_0_0_1 REGMODE_B NOREG
	 // exemplar attribute lm32_monitor_ram_0_0_1 REGMODE_A NOREG
	 // exemplar attribute lm32_monitor_ram_0_0_1 DATA_WIDTH_B 18
	 // exemplar attribute lm32_monitor_ram_0_0_1 DATA_WIDTH_A 18
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_1F 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_1E 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_1D 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_1C 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_1B 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_1A 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_19 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_18 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_17 0x0000000000000000000000000000000000000000038FF034D2038FF034C2038FF0349A038FF03EFF
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_16 0x00D00038FF034CA038FF03492038FF0348A038FF03482038FF0344A038FF03442038FF0343A038FF
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_15 0x00D6300D5A00C5803EFF0136300D0302E0803EFF02E0803EFF038FF00D5A03EFF00D630105801363
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_14 0x00D0302E0803EFF02E0803EFF038FF03EFF02E70038FF034DA0170801F100110801F100110801F10
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_13 0x0110801F100110801F100110801F100110801F100110801F100110801F100110801F100110801F08
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_12 0x02E0803EFF02E0803EFF038FF02E7802430038FF03EFF02E780110801F0803EFF030E800DE700AE7
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_11 0x00AE400AE300AE300AE300AE300AE200D0000D0000D000342000D0000D0000D000341800D0001708
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_10 0x01F100110801F100110801F100110801F100110801F100110801F0802E0803EFF0347000D0001708
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_0F 0x024700347000D00017080247002E08016E7016E4016E3016E3016E3016E3016E200DE7030E800DE7
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_0E 0x00AE703EFF010E003EFF010E003EFF010E003EFF010E0016E0016E700DE7030E800DE700AE700AE0
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_0D 0x00CE003EFF00CE003EFF00CE003EFF00CE003EFF016E700DE7030E8034700171002470030E801108
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_0C 0x01F0803470017100247000808030E80081003478011080081002478030F800AE700AE70340700AE7
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_0B 0x0344F00AE70343F00AE700AE700AE700AE600AE600AE600AE600AE500AE500AE500AE500AE400AE4
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_0A 0x00AE400AE400AE300AE300AE300AE300AE200AE200AE200AE200AE100AE100AE100AE100AE000AE0
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_09 0x00AE0030F000AE700AE70340700AE70344F00AE70343F00AE700AE700AE700AE600AE600AE600AE6
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_08 0x00AE500AE500AE500AE500AE400AE400AE400AE400AE300AE300AE300AE300AE200AE200AE200AE2
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_07 0x00AE100AE100AE100AE100AE000AE000AE0030E800DEF02EE8016E8016E800AE8016E80000800008
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_06 0x0000800008000080080800DE8016E802400016E802448016E802438016EF016EF016EF016EE016EE
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_05 0x016EE016EE016ED016ED016ED016ED016EC016EC016EC016EC016EB016EB016EB016EB016EA016EA
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_04 0x016EA016EA016E9016E9016E9016E9016E8016E8016E802600016E800DEF038FF00D0700DE702EE8
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_03 0x00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_02 0x00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_01 0x00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600
	 // exemplar attribute lm32_monitor_ram_0_1_0 INITVAL_00 0x00D000380003E0002EE0016E703E0002EE80260000D0000D0000D0000D0000D0000D0003E0002600
	 // exemplar attribute lm32_monitor_ram_0_1_0 CSDECODE_B 000
	 // exemplar attribute lm32_monitor_ram_0_1_0 CSDECODE_A 000
	 // exemplar attribute lm32_monitor_ram_0_1_0 WRITEMODE_B NORMAL
	 // exemplar attribute lm32_monitor_ram_0_1_0 WRITEMODE_A NORMAL
	 // exemplar attribute lm32_monitor_ram_0_1_0 GSR ENABLED
	 // exemplar attribute lm32_monitor_ram_0_1_0 RESETMODE ASYNC
	 // exemplar attribute lm32_monitor_ram_0_1_0 REGMODE_B NOREG
	 // exemplar attribute lm32_monitor_ram_0_1_0 REGMODE_A NOREG
	 // exemplar attribute lm32_monitor_ram_0_1_0 DATA_WIDTH_B 18
	 // exemplar attribute lm32_monitor_ram_0_1_0 DATA_WIDTH_A 18
	 // exemplar end
      end else if (lat_family == "ECP2" || lat_family == "ECP2M") begin 
	 /* Verilog netlist generated by SCUBA ispLever_v60_PROD_Build (36) */
	 /* Module Version: 3.0 */
	 /* c:\ispTOOLS6_0\ispFPGA\bin\nt\scuba.exe -w -lang verilog -synth synplify -bus_exp 7 -bb -arch ep5a00 -type bram -wp 11 -rp 1010 -addr_width 9 -data_width 32 -num_rows 512 -gsr ENABLED -writemode NORMAL -resetmode ASYNC -memfile ./rom.mem -memformat hex -e -n lm32_monitor_ram_ecp2  */
	 // synopsys translate_off
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_3F = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_3E = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_3D = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_3C = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_3B = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_3A = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_39 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_38 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_37 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_36 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_35 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_34 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_33 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_32 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_31 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_30 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_2F = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_2E = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_2D = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_2C = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_2B = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_2A = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_29 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_28 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_27 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_26 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_25 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_24 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_23 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_22 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_21 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_20 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_1F = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_1E = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_1D = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_1C = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_1B = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_1A = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_19 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_18 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_17 = 320'h00000000000000000000000000000000000000003FF8C300003FF8E300003FF90300003FF923FF5B ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_16 = 320'h1004F3FF95300003FF97300003FF99300003FF9B300003FF9D300003FF9F300003FFA1300003FFFB ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_15 = 320'h0000130001100003FF691001400000068003FF7E058003FF803FFFB300013FF7800001100001FFB3 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_14 = 320'h00000068003FF89058003FF8B3FFB93FF9B008003FFBC300000FFBE1001B000331001A0002C10019 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_13 = 320'h00035100180003510013000301001200030100110003010010000301000900030100080003010007 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_12 = 320'h010003FF97058003FFAA3FFFC00800078003FFDB3FFBD0080000004100063FFA2000000001C10004 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_11 = 320'h000083000C2001010014000183001C0000000000000001000000000000000000010000100010FFF3 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_10 = 320'h10063000481004D0003F1006D0003E1007200024100570001D10077010003FFC210000100540FFFF ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_0F = 320'h0080010000100540FFFF008000700010004000083000C2001010014000183001C0FFE40000000008 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_0E = 320'h100043FFDD100083FFDF100093FFE11000A3FFE31000B10008100040FFF8000000000C1000410008 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_0D = 320'h100083FFE7100093FFE91000A3FFEB1000B3FFED100040FFF400000200000FFFF010000000000002 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_0C = 320'h10054100000FFFF01000100FF00000100FF000000FFFE10100010000000000070300803000030090 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_0B = 320'h300003008C300003008820078100743006C2006810064000603005C2005810054000503004C20048 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_0A = 320'h10044000403003C2003810034000303002C2002810024000203001C2001810014000103000C20008 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_09 = 320'h100040000000070200802000020090200002008C20000200883007C100743006C200681006400060 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_08 = 320'h3005C2005810054000503004C2004810044000403003C2003810034000303002C200281002400020 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_07 = 320'h3001C2001810014000103000C2000810004000001F9940E000000001007410000100841000110001 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_06 = 320'h100011000110001100FF1F99410090008001008C0080010088008003007C20078000703006C20068 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_05 = 320'h10064000603005C2005810054000503004C2004810044000403003C2003810034000303002C20028 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_04 = 320'h10024000203001C2001810014000103000C200081000400000000001066C3FFC530000007F40E000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_03 = 320'h000000003B000B500800200800000A00000000000000000043000BD0080020080000120000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_02 = 320'h000000004B000C500800200800001A00000000000000000053000CD0080020080000220000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_01 = 320'h0000000081000D500800300800002A00000000000000000063000DD0080020080000320000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.INITVAL_00 = 320'h0000000091000E500800300800003A00000000000000000000000000000000000000000003F00000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.CSDECODE_B =  3'b000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.CSDECODE_A =  3'b000 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.WRITEMODE_B = "NORMAL" ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.WRITEMODE_A = "NORMAL" ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.GSR = "ENABLED" ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.RESETMODE = "ASYNC" ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.REGMODE_B = "NOREG" ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.REGMODE_A = "NOREG" ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.DATA_WIDTH_B = 18 ;
	 defparam lm32_monitor_ram_ecp2_0_0_1.DATA_WIDTH_A = 18 ;
	 // synopsys translate_on
	 DP16KB lm32_monitor_ram_ecp2_0_0_1 (.DIA0(DataInA[0]), .DIA1(DataInA[1]), 
					     .DIA2(DataInA[2]), .DIA3(DataInA[3]), .DIA4(DataInA[4]), .DIA5(DataInA[5]), 
					     .DIA6(DataInA[6]), .DIA7(DataInA[7]), .DIA8(DataInA[8]), .DIA9(DataInA[9]), 
					     .DIA10(DataInA[10]), .DIA11(DataInA[11]), .DIA12(DataInA[12]), .DIA13(DataInA[13]), 
					     .DIA14(DataInA[14]), .DIA15(DataInA[15]), .DIA16(DataInA[16]), .DIA17(DataInA[17]), 
					     .ADA0(scuba_vhi), .ADA1(scuba_vhi), .ADA2(scuba_vlo), .ADA3(scuba_vlo), 
					     .ADA4(AddressA[0]), .ADA5(AddressA[1]), .ADA6(AddressA[2]), .ADA7(AddressA[3]), 
					     .ADA8(AddressA[4]), .ADA9(AddressA[5]), .ADA10(AddressA[6]), .ADA11(AddressA[7]), 
					     .ADA12(AddressA[8]), .ADA13(scuba_vlo), .CEA(ClockEnA), .CLKA(ClockA), 
					     .WEA(WrA), .CSA0(scuba_vlo), .CSA1(scuba_vlo), .CSA2(scuba_vlo), 
					     .RSTA(ResetA), .DIB0(DataInB[0]), .DIB1(DataInB[1]), .DIB2(DataInB[2]), 
					     .DIB3(DataInB[3]), .DIB4(DataInB[4]), .DIB5(DataInB[5]), .DIB6(DataInB[6]), 
					     .DIB7(DataInB[7]), .DIB8(DataInB[8]), .DIB9(DataInB[9]), .DIB10(DataInB[10]), 
					     .DIB11(DataInB[11]), .DIB12(DataInB[12]), .DIB13(DataInB[13]), .DIB14(DataInB[14]), 
					     .DIB15(DataInB[15]), .DIB16(DataInB[16]), .DIB17(DataInB[17]), .ADB0(scuba_vhi), 
					     .ADB1(scuba_vhi), .ADB2(scuba_vlo), .ADB3(scuba_vlo), .ADB4(AddressB[0]), 
					     .ADB5(AddressB[1]), .ADB6(AddressB[2]), .ADB7(AddressB[3]), .ADB8(AddressB[4]), 
					     .ADB9(AddressB[5]), .ADB10(AddressB[6]), .ADB11(AddressB[7]), .ADB12(AddressB[8]), 
					     .ADB13(scuba_vlo), .CEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB0(scuba_vlo), 
					     .CSB1(scuba_vlo), .CSB2(scuba_vlo), .RSTB(ResetB), .DOA0(QA[0]), 
					     .DOA1(QA[1]), .DOA2(QA[2]), .DOA3(QA[3]), .DOA4(QA[4]), .DOA5(QA[5]), 
					     .DOA6(QA[6]), .DOA7(QA[7]), .DOA8(QA[8]), .DOA9(QA[9]), .DOA10(QA[10]), 
					     .DOA11(QA[11]), .DOA12(QA[12]), .DOA13(QA[13]), .DOA14(QA[14]), 
					     .DOA15(QA[15]), .DOA16(QA[16]), .DOA17(QA[17]), .DOB0(QB[0]), .DOB1(QB[1]), 
					     .DOB2(QB[2]), .DOB3(QB[3]), .DOB4(QB[4]), .DOB5(QB[5]), .DOB6(QB[6]), 
					     .DOB7(QB[7]), .DOB8(QB[8]), .DOB9(QB[9]), .DOB10(QB[10]), .DOB11(QB[11]), 
					     .DOB12(QB[12]), .DOB13(QB[13]), .DOB14(QB[14]), .DOB15(QB[15]), 
					     .DOB16(QB[16]), .DOB17(QB[17]))
           /* synthesis MEM_LPC_FILE="lm32_monitor_ram_ecp2.lpc" */
           /* synthesis MEM_INIT_FILE="rom.mem" */
           /* synthesis INITVAL_3F="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_3E="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_3D="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_3C="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_3B="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_3A="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_39="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_38="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_37="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_36="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_35="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_34="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_33="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_32="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_31="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_30="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2F="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2E="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2D="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2C="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2B="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2A="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_29="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_28="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_27="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_26="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_25="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_24="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_23="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_22="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_21="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_20="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1F="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1E="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1D="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1C="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1B="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1A="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_19="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_18="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_17="0x00000000000000000000000000000000000000003FF8C300003FF8E300003FF90300003FF923FF5B" */
           /* synthesis INITVAL_16="0x1004F3FF95300003FF97300003FF99300003FF9B300003FF9D300003FF9F300003FFA1300003FFFB" */
           /* synthesis INITVAL_15="0x0000130001100003FF691001400000068003FF7E058003FF803FFFB300013FF7800001100001FFB3" */
           /* synthesis INITVAL_14="0x00000068003FF89058003FF8B3FFB93FF9B008003FFBC300000FFBE1001B000331001A0002C10019" */
           /* synthesis INITVAL_13="0x00035100180003510013000301001200030100110003010010000301000900030100080003010007" */
           /* synthesis INITVAL_12="0x010003FF97058003FFAA3FFFC00800078003FFDB3FFBD0080000004100063FFA2000000001C10004" */
           /* synthesis INITVAL_11="0x000083000C2001010014000183001C0000000000000001000000000000000000010000100010FFF3" */
           /* synthesis INITVAL_10="0x10063000481004D0003F1006D0003E1007200024100570001D10077010003FFC210000100540FFFF" */
           /* synthesis INITVAL_0F="0x0080010000100540FFFF008000700010004000083000C2001010014000183001C0FFE40000000008" */
           /* synthesis INITVAL_0E="0x100043FFDD100083FFDF100093FFE11000A3FFE31000B10008100040FFF8000000000C1000410008" */
           /* synthesis INITVAL_0D="0x100083FFE7100093FFE91000A3FFEB1000B3FFED100040FFF400000200000FFFF010000000000002" */
           /* synthesis INITVAL_0C="0x10054100000FFFF01000100FF00000100FF000000FFFE10100010000000000070300803000030090" */
           /* synthesis INITVAL_0B="0x300003008C300003008820078100743006C2006810064000603005C2005810054000503004C20048" */
           /* synthesis INITVAL_0A="0x10044000403003C2003810034000303002C2002810024000203001C2001810014000103000C20008" */
           /* synthesis INITVAL_09="0x100040000000070200802000020090200002008C20000200883007C100743006C200681006400060" */
           /* synthesis INITVAL_08="0x3005C2005810054000503004C2004810044000403003C2003810034000303002C200281002400020" */
           /* synthesis INITVAL_07="0x3001C2001810014000103000C2000810004000001F9940E000000001007410000100841000110001" */
           /* synthesis INITVAL_06="0x100011000110001100FF1F99410090008001008C0080010088008003007C20078000703006C20068" */
           /* synthesis INITVAL_05="0x10064000603005C2005810054000503004C2004810044000403003C2003810034000303002C20028" */
           /* synthesis INITVAL_04="0x10024000203001C2001810014000103000C200081000400000000001066C3FFC530000007F40E000" */
           /* synthesis INITVAL_03="0x000000003B000B500800200800000A00000000000000000043000BD0080020080000120000000000" */
           /* synthesis INITVAL_02="0x000000004B000C500800200800001A00000000000000000053000CD0080020080000220000000000" */
           /* synthesis INITVAL_01="0x0000000081000D500800300800002A00000000000000000063000DD0080020080000320000000000" */
           /* synthesis INITVAL_00="0x0000000091000E500800300800003A00000000000000000000000000000000000000000003F00000" */
           /* synthesis CSDECODE_B="0b000" */
           /* synthesis CSDECODE_A="0b000" */
           /* synthesis WRITEMODE_B="NORMAL" */
           /* synthesis WRITEMODE_A="NORMAL" */
           /* synthesis GSR="ENABLED" */
           /* synthesis RESETMODE="ASYNC" */
           /* synthesis REGMODE_B="NOREG" */
           /* synthesis REGMODE_A="NOREG" */
           /* synthesis DATA_WIDTH_B="18" */
           /* synthesis DATA_WIDTH_A="18" */;

	 VHI scuba_vhi_inst (.Z(scuba_vhi));

	 VLO scuba_vlo_inst (.Z(scuba_vlo));

	 // synopsys translate_off
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_3F = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_3E = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_3D = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_3C = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_3B = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_3A = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_39 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_38 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_37 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_36 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_35 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_34 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_33 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_32 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_31 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_30 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_2F = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_2E = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_2D = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_2C = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_2B = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_2A = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_29 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_28 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_27 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_26 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_25 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_24 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_23 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_22 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_21 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_20 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_1F = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_1E = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_1D = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_1C = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_1B = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_1A = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_19 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_18 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_17 = 320'h0000000000000000000000000000000000000000038FF034D2038FF034C2038FF0349A038FF03EFF ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_16 = 320'h00D00038FF034CA038FF03492038FF0348A038FF03482038FF0344A038FF03442038FF0343A038FF ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_15 = 320'h00D6300D5A00C5803EFF0136300D0302E0803EFF02E0803EFF038FF00D5A03EFF00D630105801363 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_14 = 320'h00D0302E0803EFF02E0803EFF038FF03EFF02E70038FF034DA0170801F100110801F100110801F10 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_13 = 320'h0110801F100110801F100110801F100110801F100110801F100110801F100110801F100110801F08 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_12 = 320'h02E0803EFF02E0803EFF038FF02E7802430038FF03EFF02E780110801F0803EFF030E800DE700AE7 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_11 = 320'h00AE400AE300AE300AE300AE300AE200D0000D0000D000342000D0000D0000D000341800D0001708 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_10 = 320'h01F100110801F100110801F100110801F100110801F100110801F0802E0803EFF0347000D0001708 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_0F = 320'h024700347000D00017080247002E08016E7016E4016E3016E3016E3016E3016E200DE7030E800DE7 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_0E = 320'h00AE703EFF010E003EFF010E003EFF010E003EFF010E0016E0016E700DE7030E800DE700AE700AE0 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_0D = 320'h00CE003EFF00CE003EFF00CE003EFF00CE003EFF016E700DE7030E8034700171002470030E801108 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_0C = 320'h01F0803470017100247000808030E80081003478011080081002478030F800AE700AE70340700AE7 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_0B = 320'h0344F00AE70343F00AE700AE700AE700AE600AE600AE600AE600AE500AE500AE500AE500AE400AE4 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_0A = 320'h00AE400AE400AE300AE300AE300AE300AE200AE200AE200AE200AE100AE100AE100AE100AE000AE0 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_09 = 320'h00AE0030F000AE700AE70340700AE70344F00AE70343F00AE700AE700AE700AE600AE600AE600AE6 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_08 = 320'h00AE500AE500AE500AE500AE400AE400AE400AE400AE300AE300AE300AE300AE200AE200AE200AE2 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_07 = 320'h00AE100AE100AE100AE100AE000AE000AE0030E800DEF02EE8016E8016E800AE8016E80000800008 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_06 = 320'h0000800008000080080800DE8016E802400016E802448016E802438016EF016EF016EF016EE016EE ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_05 = 320'h016EE016EE016ED016ED016ED016ED016EC016EC016EC016EC016EB016EB016EB016EB016EA016EA ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_04 = 320'h016EA016EA016E9016E9016E9016E9016E8016E8016E802600016E800DEF038FF00D0700DE702EE8 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_03 = 320'h00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_02 = 320'h00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_01 = 320'h00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.INITVAL_00 = 320'h00D000380003E0002EE0016E703E0002EE80260000D0000D0000D0000D0000D0000D0003E0002600 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.CSDECODE_B =  3'b000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.CSDECODE_A =  3'b000 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.WRITEMODE_B = "NORMAL" ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.WRITEMODE_A = "NORMAL" ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.GSR = "ENABLED" ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.RESETMODE = "ASYNC" ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.REGMODE_B = "NOREG" ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.REGMODE_A = "NOREG" ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.DATA_WIDTH_B = 18 ;
	 defparam lm32_monitor_ram_ecp2_0_1_0.DATA_WIDTH_A = 18 ;
	 // synopsys translate_on
	 DP16KB lm32_monitor_ram_ecp2_0_1_0 (.DIA0(DataInA[18]), .DIA1(DataInA[19]), 
					     .DIA2(DataInA[20]), .DIA3(DataInA[21]), .DIA4(DataInA[22]), .DIA5(DataInA[23]), 
					     .DIA6(DataInA[24]), .DIA7(DataInA[25]), .DIA8(DataInA[26]), .DIA9(DataInA[27]), 
					     .DIA10(DataInA[28]), .DIA11(DataInA[29]), .DIA12(DataInA[30]), .DIA13(DataInA[31]), 
					     .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), .DIA17(scuba_vlo), 
					     .ADA0(scuba_vhi), .ADA1(scuba_vhi), .ADA2(scuba_vlo), .ADA3(scuba_vlo), 
					     .ADA4(AddressA[0]), .ADA5(AddressA[1]), .ADA6(AddressA[2]), .ADA7(AddressA[3]), 
					     .ADA8(AddressA[4]), .ADA9(AddressA[5]), .ADA10(AddressA[6]), .ADA11(AddressA[7]), 
					     .ADA12(AddressA[8]), .ADA13(scuba_vlo), .CEA(ClockEnA), .CLKA(ClockA), 
					     .WEA(WrA), .CSA0(scuba_vlo), .CSA1(scuba_vlo), .CSA2(scuba_vlo), 
					     .RSTA(ResetA), .DIB0(DataInB[18]), .DIB1(DataInB[19]), .DIB2(DataInB[20]), 
					     .DIB3(DataInB[21]), .DIB4(DataInB[22]), .DIB5(DataInB[23]), .DIB6(DataInB[24]), 
					     .DIB7(DataInB[25]), .DIB8(DataInB[26]), .DIB9(DataInB[27]), .DIB10(DataInB[28]), 
					     .DIB11(DataInB[29]), .DIB12(DataInB[30]), .DIB13(DataInB[31]), .DIB14(scuba_vlo), 
					     .DIB15(scuba_vlo), .DIB16(scuba_vlo), .DIB17(scuba_vlo), .ADB0(scuba_vhi), 
					     .ADB1(scuba_vhi), .ADB2(scuba_vlo), .ADB3(scuba_vlo), .ADB4(AddressB[0]), 
					     .ADB5(AddressB[1]), .ADB6(AddressB[2]), .ADB7(AddressB[3]), .ADB8(AddressB[4]), 
					     .ADB9(AddressB[5]), .ADB10(AddressB[6]), .ADB11(AddressB[7]), .ADB12(AddressB[8]), 
					     .ADB13(scuba_vlo), .CEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB0(scuba_vlo), 
					     .CSB1(scuba_vlo), .CSB2(scuba_vlo), .RSTB(ResetB), .DOA0(QA[18]), 
					     .DOA1(QA[19]), .DOA2(QA[20]), .DOA3(QA[21]), .DOA4(QA[22]), .DOA5(QA[23]), 
					     .DOA6(QA[24]), .DOA7(QA[25]), .DOA8(QA[26]), .DOA9(QA[27]), .DOA10(QA[28]), 
					     .DOA11(QA[29]), .DOA12(QA[30]), .DOA13(QA[31]), .DOA14(), .DOA15(), 
					     .DOA16(), .DOA17(), .DOB0(QB[18]), .DOB1(QB[19]), .DOB2(QB[20]), 
					     .DOB3(QB[21]), .DOB4(QB[22]), .DOB5(QB[23]), .DOB6(QB[24]), .DOB7(QB[25]), 
					     .DOB8(QB[26]), .DOB9(QB[27]), .DOB10(QB[28]), .DOB11(QB[29]), .DOB12(QB[30]), 
					     .DOB13(QB[31]), .DOB14(), .DOB15(), .DOB16(), .DOB17())
           /* synthesis MEM_LPC_FILE="lm32_monitor_ram_ecp2.lpc" */
           /* synthesis MEM_INIT_FILE="rom.mem" */
           /* synthesis INITVAL_3F="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_3E="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_3D="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_3C="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_3B="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_3A="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_39="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_38="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_37="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_36="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_35="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_34="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_33="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_32="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_31="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_30="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2F="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2E="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2D="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2C="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2B="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2A="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_29="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_28="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_27="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_26="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_25="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_24="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_23="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_22="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_21="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_20="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1F="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1E="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1D="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1C="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1B="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1A="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_19="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_18="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_17="0x0000000000000000000000000000000000000000038FF034D2038FF034C2038FF0349A038FF03EFF" */
           /* synthesis INITVAL_16="0x00D00038FF034CA038FF03492038FF0348A038FF03482038FF0344A038FF03442038FF0343A038FF" */
           /* synthesis INITVAL_15="0x00D6300D5A00C5803EFF0136300D0302E0803EFF02E0803EFF038FF00D5A03EFF00D630105801363" */
           /* synthesis INITVAL_14="0x00D0302E0803EFF02E0803EFF038FF03EFF02E70038FF034DA0170801F100110801F100110801F10" */
           /* synthesis INITVAL_13="0x0110801F100110801F100110801F100110801F100110801F100110801F100110801F100110801F08" */
           /* synthesis INITVAL_12="0x02E0803EFF02E0803EFF038FF02E7802430038FF03EFF02E780110801F0803EFF030E800DE700AE7" */
           /* synthesis INITVAL_11="0x00AE400AE300AE300AE300AE300AE200D0000D0000D000342000D0000D0000D000341800D0001708" */
           /* synthesis INITVAL_10="0x01F100110801F100110801F100110801F100110801F100110801F0802E0803EFF0347000D0001708" */
           /* synthesis INITVAL_0F="0x024700347000D00017080247002E08016E7016E4016E3016E3016E3016E3016E200DE7030E800DE7" */
           /* synthesis INITVAL_0E="0x00AE703EFF010E003EFF010E003EFF010E003EFF010E0016E0016E700DE7030E800DE700AE700AE0" */
           /* synthesis INITVAL_0D="0x00CE003EFF00CE003EFF00CE003EFF00CE003EFF016E700DE7030E8034700171002470030E801108" */
           /* synthesis INITVAL_0C="0x01F0803470017100247000808030E80081003478011080081002478030F800AE700AE70340700AE7" */
           /* synthesis INITVAL_0B="0x0344F00AE70343F00AE700AE700AE700AE600AE600AE600AE600AE500AE500AE500AE500AE400AE4" */
           /* synthesis INITVAL_0A="0x00AE400AE400AE300AE300AE300AE300AE200AE200AE200AE200AE100AE100AE100AE100AE000AE0" */
           /* synthesis INITVAL_09="0x00AE0030F000AE700AE70340700AE70344F00AE70343F00AE700AE700AE700AE600AE600AE600AE6" */
           /* synthesis INITVAL_08="0x00AE500AE500AE500AE500AE400AE400AE400AE400AE300AE300AE300AE300AE200AE200AE200AE2" */
           /* synthesis INITVAL_07="0x00AE100AE100AE100AE100AE000AE000AE0030E800DEF02EE8016E8016E800AE8016E80000800008" */
           /* synthesis INITVAL_06="0x0000800008000080080800DE8016E802400016E802448016E802438016EF016EF016EF016EE016EE" */
           /* synthesis INITVAL_05="0x016EE016EE016ED016ED016ED016ED016EC016EC016EC016EC016EB016EB016EB016EB016EA016EA" */
           /* synthesis INITVAL_04="0x016EA016EA016E9016E9016E9016E9016E8016E8016E802600016E800DEF038FF00D0700DE702EE8" */
           /* synthesis INITVAL_03="0x00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600" */
           /* synthesis INITVAL_02="0x00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600" */
           /* synthesis INITVAL_01="0x00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600" */
           /* synthesis INITVAL_00="0x00D000380003E0002EE0016E703E0002EE80260000D0000D0000D0000D0000D0000D0003E0002600" */
           /* synthesis CSDECODE_B="0b000" */
           /* synthesis CSDECODE_A="0b000" */
           /* synthesis WRITEMODE_B="NORMAL" */
           /* synthesis WRITEMODE_A="NORMAL" */
           /* synthesis GSR="ENABLED" */
           /* synthesis RESETMODE="ASYNC" */
           /* synthesis REGMODE_B="NOREG" */
           /* synthesis REGMODE_A="NOREG" */
           /* synthesis DATA_WIDTH_B="18" */
           /* synthesis DATA_WIDTH_A="18" */;



	 // exemplar begin
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 MEM_LPC_FILE lm32_monitor_ram_ecp2.lpc
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 MEM_INIT_FILE rom.mem
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_3F 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_3E 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_3D 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_3C 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_3B 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_3A 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_39 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_38 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_37 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_36 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_35 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_34 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_33 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_32 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_31 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_30 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_2F 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_2E 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_2D 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_2C 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_2B 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_2A 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_29 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_28 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_27 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_26 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_25 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_24 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_23 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_22 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_21 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_20 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_1F 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_1E 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_1D 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_1C 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_1B 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_1A 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_19 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_18 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_17 0x00000000000000000000000000000000000000003FF8C300003FF8E300003FF90300003FF923FF5B
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_16 0x1004F3FF95300003FF97300003FF99300003FF9B300003FF9D300003FF9F300003FFA1300003FFFB
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_15 0x0000130001100003FF691001400000068003FF7E058003FF803FFFB300013FF7800001100001FFB3
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_14 0x00000068003FF89058003FF8B3FFB93FF9B008003FFBC300000FFBE1001B000331001A0002C10019
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_13 0x00035100180003510013000301001200030100110003010010000301000900030100080003010007
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_12 0x010003FF97058003FFAA3FFFC00800078003FFDB3FFBD0080000004100063FFA2000000001C10004
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_11 0x000083000C2001010014000183001C0000000000000001000000000000000000010000100010FFF3
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_10 0x10063000481004D0003F1006D0003E1007200024100570001D10077010003FFC210000100540FFFF
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_0F 0x0080010000100540FFFF008000700010004000083000C2001010014000183001C0FFE40000000008
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_0E 0x100043FFDD100083FFDF100093FFE11000A3FFE31000B10008100040FFF8000000000C1000410008
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_0D 0x100083FFE7100093FFE91000A3FFEB1000B3FFED100040FFF400000200000FFFF010000000000002
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_0C 0x10054100000FFFF01000100FF00000100FF000000FFFE10100010000000000070300803000030090
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_0B 0x300003008C300003008820078100743006C2006810064000603005C2005810054000503004C20048
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_0A 0x10044000403003C2003810034000303002C2002810024000203001C2001810014000103000C20008
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_09 0x100040000000070200802000020090200002008C20000200883007C100743006C200681006400060
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_08 0x3005C2005810054000503004C2004810044000403003C2003810034000303002C200281002400020
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_07 0x3001C2001810014000103000C2000810004000001F9940E000000001007410000100841000110001
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_06 0x100011000110001100FF1F99410090008001008C0080010088008003007C20078000703006C20068
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_05 0x10064000603005C2005810054000503004C2004810044000403003C2003810034000303002C20028
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_04 0x10024000203001C2001810014000103000C200081000400000000001066C3FFC530000007F40E000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_03 0x000000003B000B500800200800000A00000000000000000043000BD0080020080000120000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_02 0x000000004B000C500800200800001A00000000000000000053000CD0080020080000220000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_01 0x0000000081000D500800300800002A00000000000000000063000DD0080020080000320000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 INITVAL_00 0x0000000091000E500800300800003A00000000000000000000000000000000000000000003F00000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 CSDECODE_B 0b000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 CSDECODE_A 0b000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 WRITEMODE_B NORMAL
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 WRITEMODE_A NORMAL
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 GSR ENABLED
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 RESETMODE ASYNC
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 REGMODE_B NOREG
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 REGMODE_A NOREG
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 DATA_WIDTH_B 18
	 // exemplar attribute lm32_monitor_ram_ecp2_0_0_1 DATA_WIDTH_A 18
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 MEM_LPC_FILE lm32_monitor_ram_ecp2.lpc
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 MEM_INIT_FILE rom.mem
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_3F 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_3E 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_3D 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_3C 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_3B 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_3A 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_39 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_38 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_37 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_36 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_35 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_34 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_33 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_32 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_31 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_30 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_2F 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_2E 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_2D 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_2C 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_2B 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_2A 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_29 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_28 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_27 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_26 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_25 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_24 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_23 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_22 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_21 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_20 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_1F 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_1E 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_1D 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_1C 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_1B 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_1A 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_19 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_18 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_17 0x0000000000000000000000000000000000000000038FF034D2038FF034C2038FF0349A038FF03EFF
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_16 0x00D00038FF034CA038FF03492038FF0348A038FF03482038FF0344A038FF03442038FF0343A038FF
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_15 0x00D6300D5A00C5803EFF0136300D0302E0803EFF02E0803EFF038FF00D5A03EFF00D630105801363
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_14 0x00D0302E0803EFF02E0803EFF038FF03EFF02E70038FF034DA0170801F100110801F100110801F10
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_13 0x0110801F100110801F100110801F100110801F100110801F100110801F100110801F100110801F08
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_12 0x02E0803EFF02E0803EFF038FF02E7802430038FF03EFF02E780110801F0803EFF030E800DE700AE7
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_11 0x00AE400AE300AE300AE300AE300AE200D0000D0000D000342000D0000D0000D000341800D0001708
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_10 0x01F100110801F100110801F100110801F100110801F100110801F0802E0803EFF0347000D0001708
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_0F 0x024700347000D00017080247002E08016E7016E4016E3016E3016E3016E3016E200DE7030E800DE7
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_0E 0x00AE703EFF010E003EFF010E003EFF010E003EFF010E0016E0016E700DE7030E800DE700AE700AE0
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_0D 0x00CE003EFF00CE003EFF00CE003EFF00CE003EFF016E700DE7030E8034700171002470030E801108
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_0C 0x01F0803470017100247000808030E80081003478011080081002478030F800AE700AE70340700AE7
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_0B 0x0344F00AE70343F00AE700AE700AE700AE600AE600AE600AE600AE500AE500AE500AE500AE400AE4
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_0A 0x00AE400AE400AE300AE300AE300AE300AE200AE200AE200AE200AE100AE100AE100AE100AE000AE0
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_09 0x00AE0030F000AE700AE70340700AE70344F00AE70343F00AE700AE700AE700AE600AE600AE600AE6
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_08 0x00AE500AE500AE500AE500AE400AE400AE400AE400AE300AE300AE300AE300AE200AE200AE200AE2
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_07 0x00AE100AE100AE100AE100AE000AE000AE0030E800DEF02EE8016E8016E800AE8016E80000800008
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_06 0x0000800008000080080800DE8016E802400016E802448016E802438016EF016EF016EF016EE016EE
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_05 0x016EE016EE016ED016ED016ED016ED016EC016EC016EC016EC016EB016EB016EB016EB016EA016EA
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_04 0x016EA016EA016E9016E9016E9016E9016E8016E8016E802600016E800DEF038FF00D0700DE702EE8
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_03 0x00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_02 0x00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_01 0x00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 INITVAL_00 0x00D000380003E0002EE0016E703E0002EE80260000D0000D0000D0000D0000D0000D0003E0002600
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 CSDECODE_B 0b000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 CSDECODE_A 0b000
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 WRITEMODE_B NORMAL
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 WRITEMODE_A NORMAL
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 GSR ENABLED
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 RESETMODE ASYNC
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 REGMODE_B NOREG
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 REGMODE_A NOREG
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 DATA_WIDTH_B 18
	 // exemplar attribute lm32_monitor_ram_ecp2_0_1_0 DATA_WIDTH_A 18
	 // exemplar end
      end   else if (lat_family == "SC" || lat_family == "SCM") begin 
	 // synopsys translate_off
	 defparam sc_rom_monitor_0_0_1.INITVAL_3F = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_3E = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_3D = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_3C = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_3B = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_3A = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_39 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_38 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_37 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_36 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_35 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_34 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_33 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_32 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_31 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_30 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_2F = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_2E = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_2D = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_2C = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_2B = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_2A = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_29 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_28 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_27 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_26 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_25 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_24 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_23 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_22 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_21 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_20 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_1F = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_1E = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_1D = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_1C = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_1B = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_1A = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_19 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_18 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_17 = 320'h00000000000000000000000000000000000000003FF8C300003FF8E300003FF90300003FF923FF5B ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_16 = 320'h1004F3FF95300003FF97300003FF99300003FF9B300003FF9D300003FF9F300003FFA1300003FFFB ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_15 = 320'h0000130001100003FF691001400000068003FF7E058003FF803FFFB300013FF7800001100001FFB3 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_14 = 320'h00000068003FF89058003FF8B3FFB93FF9B008003FFBC300000FFBE1001B000331001A0002C10019 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_13 = 320'h00035100180003510013000301001200030100110003010010000301000900030100080003010007 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_12 = 320'h010003FF97058003FFAA3FFFC00800078003FFDB3FFBD0080000004100063FFA2000000001C10004 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_11 = 320'h000083000C2001010014000183001C0000000000000001000000000000000000010000100010FFF3 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_10 = 320'h10063000481004D0003F1006D0003E1007200024100570001D10077010003FFC210000100540FFFF ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_0F = 320'h0080010000100540FFFF008000700010004000083000C2001010014000183001C0FFE40000000008 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_0E = 320'h100043FFDD100083FFDF100093FFE11000A3FFE31000B10008100040FFF8000000000C1000410008 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_0D = 320'h100083FFE7100093FFE91000A3FFEB1000B3FFED100040FFF400000200000FFFF010000000000002 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_0C = 320'h10054100000FFFF01000100FF00000100FF000000FFFE10100010000000000070300803000030090 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_0B = 320'h300003008C300003008820078100743006C2006810064000603005C2005810054000503004C20048 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_0A = 320'h10044000403003C2003810034000303002C2002810024000203001C2001810014000103000C20008 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_09 = 320'h100040000000070200802000020090200002008C20000200883007C100743006C200681006400060 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_08 = 320'h3005C2005810054000503004C2004810044000403003C2003810034000303002C200281002400020 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_07 = 320'h3001C2001810014000103000C2000810004000001F9940E000000001007410000100841000110001 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_06 = 320'h100011000110001100FF1F99410090008001008C0080010088008003007C20078000703006C20068 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_05 = 320'h10064000603005C2005810054000503004C2004810044000403003C2003810034000303002C20028 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_04 = 320'h10024000203001C2001810014000103000C200081000400000000001066C3FFC530000007F40E000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_03 = 320'h000000003B000B500800200800000A00000000000000000043000BD0080020080000120000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_02 = 320'h000000004B000C500800200800001A00000000000000000053000CD0080020080000220000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_01 = 320'h0000000081000D500800300800002A00000000000000000063000DD0080020080000320000000000 ;
	 defparam sc_rom_monitor_0_0_1.INITVAL_00 = 320'h0000000091000E500800300800003A00000000000000000000000000000000000000000003F00000 ;
	 defparam sc_rom_monitor_0_0_1.CSDECODE_B =  3'b000 ;
	 defparam sc_rom_monitor_0_0_1.CSDECODE_A =  3'b000 ;
	 defparam sc_rom_monitor_0_0_1.WRITEMODE_B = "NORMAL" ;
	 defparam sc_rom_monitor_0_0_1.WRITEMODE_A = "NORMAL" ;
	 defparam sc_rom_monitor_0_0_1.GSR = "ENABLED" ;
	 defparam sc_rom_monitor_0_0_1.RESETMODE = "ASYNC" ;
	 defparam sc_rom_monitor_0_0_1.REGMODE_B = "NOREG" ;
	 defparam sc_rom_monitor_0_0_1.REGMODE_A = "NOREG" ;
	 defparam sc_rom_monitor_0_0_1.DATA_WIDTH_B = 18 ;
	 defparam sc_rom_monitor_0_0_1.DATA_WIDTH_A = 18 ;
	 // synopsys translate_on
	 DP16KA sc_rom_monitor_0_0_1 (.DIA0(DataInA[0]), .DIA1(DataInA[1]), .DIA2(DataInA[2]), 
				      .DIA3(DataInA[3]), .DIA4(DataInA[4]), .DIA5(DataInA[5]), .DIA6(DataInA[6]), 
				      .DIA7(DataInA[7]), .DIA8(DataInA[8]), .DIA9(DataInA[9]), .DIA10(DataInA[10]), 
				      .DIA11(DataInA[11]), .DIA12(DataInA[12]), .DIA13(DataInA[13]), .DIA14(DataInA[14]), 
				      .DIA15(DataInA[15]), .DIA16(DataInA[16]), .DIA17(DataInA[17]), .ADA0(scuba_vhi), 
				      .ADA1(scuba_vhi), .ADA2(scuba_vlo), .ADA3(scuba_vlo), .ADA4(AddressA[0]), 
				      .ADA5(AddressA[1]), .ADA6(AddressA[2]), .ADA7(AddressA[3]), .ADA8(AddressA[4]), 
				      .ADA9(AddressA[5]), .ADA10(AddressA[6]), .ADA11(AddressA[7]), .ADA12(AddressA[8]), 
				      .ADA13(scuba_vlo), .CEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA0(scuba_vlo), 
				      .CSA1(scuba_vlo), .CSA2(scuba_vlo), .RSTA(ResetA), .DIB0(DataInB[0]), 
				      .DIB1(DataInB[1]), .DIB2(DataInB[2]), .DIB3(DataInB[3]), .DIB4(DataInB[4]), 
				      .DIB5(DataInB[5]), .DIB6(DataInB[6]), .DIB7(DataInB[7]), .DIB8(DataInB[8]), 
				      .DIB9(DataInB[9]), .DIB10(DataInB[10]), .DIB11(DataInB[11]), .DIB12(DataInB[12]), 
				      .DIB13(DataInB[13]), .DIB14(DataInB[14]), .DIB15(DataInB[15]), .DIB16(DataInB[16]), 
				      .DIB17(DataInB[17]), .ADB0(scuba_vhi), .ADB1(scuba_vhi), .ADB2(scuba_vlo), 
				      .ADB3(scuba_vlo), .ADB4(AddressB[0]), .ADB5(AddressB[1]), .ADB6(AddressB[2]), 
				      .ADB7(AddressB[3]), .ADB8(AddressB[4]), .ADB9(AddressB[5]), .ADB10(AddressB[6]), 
				      .ADB11(AddressB[7]), .ADB12(AddressB[8]), .ADB13(scuba_vlo), .CEB(ClockEnB), 
				      .CLKB(ClockB), .WEB(WrB), .CSB0(scuba_vlo), .CSB1(scuba_vlo), .CSB2(scuba_vlo), 
				      .RSTB(ResetB), .DOA0(QA[0]), .DOA1(QA[1]), .DOA2(QA[2]), .DOA3(QA[3]), 
				      .DOA4(QA[4]), .DOA5(QA[5]), .DOA6(QA[6]), .DOA7(QA[7]), .DOA8(QA[8]), 
				      .DOA9(QA[9]), .DOA10(QA[10]), .DOA11(QA[11]), .DOA12(QA[12]), .DOA13(QA[13]), 
				      .DOA14(QA[14]), .DOA15(QA[15]), .DOA16(QA[16]), .DOA17(QA[17]), 
				      .DOB0(QB[0]), .DOB1(QB[1]), .DOB2(QB[2]), .DOB3(QB[3]), .DOB4(QB[4]), 
				      .DOB5(QB[5]), .DOB6(QB[6]), .DOB7(QB[7]), .DOB8(QB[8]), .DOB9(QB[9]), 
				      .DOB10(QB[10]), .DOB11(QB[11]), .DOB12(QB[12]), .DOB13(QB[13]), 
				      .DOB14(QB[14]), .DOB15(QB[15]), .DOB16(QB[16]), .DOB17(QB[17]))
           /* synthesis MEM_LPC_FILE="sc_rom_monitor.lpc" */
           /* synthesis MEM_INIT_FILE="rom.mem" */
           /* synthesis INITVAL_3F="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_3E="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_3D="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_3C="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_3B="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_3A="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_39="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_38="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_37="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_36="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_35="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_34="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_33="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_32="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_31="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_30="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2F="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2E="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2D="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2C="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2B="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2A="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_29="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_28="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_27="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_26="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_25="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_24="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_23="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_22="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_21="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_20="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1F="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1E="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1D="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1C="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1B="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1A="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_19="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_18="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_17="0x00000000000000000000000000000000000000003FF8C300003FF8E300003FF90300003FF923FF5B" */
           /* synthesis INITVAL_16="0x1004F3FF95300003FF97300003FF99300003FF9B300003FF9D300003FF9F300003FFA1300003FFFB" */
           /* synthesis INITVAL_15="0x0000130001100003FF691001400000068003FF7E058003FF803FFFB300013FF7800001100001FFB3" */
           /* synthesis INITVAL_14="0x00000068003FF89058003FF8B3FFB93FF9B008003FFBC300000FFBE1001B000331001A0002C10019" */
           /* synthesis INITVAL_13="0x00035100180003510013000301001200030100110003010010000301000900030100080003010007" */
           /* synthesis INITVAL_12="0x010003FF97058003FFAA3FFFC00800078003FFDB3FFBD0080000004100063FFA2000000001C10004" */
           /* synthesis INITVAL_11="0x000083000C2001010014000183001C0000000000000001000000000000000000010000100010FFF3" */
           /* synthesis INITVAL_10="0x10063000481004D0003F1006D0003E1007200024100570001D10077010003FFC210000100540FFFF" */
           /* synthesis INITVAL_0F="0x0080010000100540FFFF008000700010004000083000C2001010014000183001C0FFE40000000008" */
           /* synthesis INITVAL_0E="0x100043FFDD100083FFDF100093FFE11000A3FFE31000B10008100040FFF8000000000C1000410008" */
           /* synthesis INITVAL_0D="0x100083FFE7100093FFE91000A3FFEB1000B3FFED100040FFF400000200000FFFF010000000000002" */
           /* synthesis INITVAL_0C="0x10054100000FFFF01000100FF00000100FF000000FFFE10100010000000000070300803000030090" */
           /* synthesis INITVAL_0B="0x300003008C300003008820078100743006C2006810064000603005C2005810054000503004C20048" */
           /* synthesis INITVAL_0A="0x10044000403003C2003810034000303002C2002810024000203001C2001810014000103000C20008" */
           /* synthesis INITVAL_09="0x100040000000070200802000020090200002008C20000200883007C100743006C200681006400060" */
           /* synthesis INITVAL_08="0x3005C2005810054000503004C2004810044000403003C2003810034000303002C200281002400020" */
           /* synthesis INITVAL_07="0x3001C2001810014000103000C2000810004000001F9940E000000001007410000100841000110001" */
           /* synthesis INITVAL_06="0x100011000110001100FF1F99410090008001008C0080010088008003007C20078000703006C20068" */
           /* synthesis INITVAL_05="0x10064000603005C2005810054000503004C2004810044000403003C2003810034000303002C20028" */
           /* synthesis INITVAL_04="0x10024000203001C2001810014000103000C200081000400000000001066C3FFC530000007F40E000" */
           /* synthesis INITVAL_03="0x000000003B000B500800200800000A00000000000000000043000BD0080020080000120000000000" */
           /* synthesis INITVAL_02="0x000000004B000C500800200800001A00000000000000000053000CD0080020080000220000000000" */
           /* synthesis INITVAL_01="0x0000000081000D500800300800002A00000000000000000063000DD0080020080000320000000000" */
           /* synthesis INITVAL_00="0x0000000091000E500800300800003A00000000000000000000000000000000000000000003F00000" */
           /* synthesis CSDECODE_B="0b000" */
           /* synthesis CSDECODE_A="0b000" */
           /* synthesis WRITEMODE_B="NORMAL" */
           /* synthesis WRITEMODE_A="NORMAL" */
           /* synthesis GSR="ENABLED" */
           /* synthesis RESETMODE="ASYNC" */
           /* synthesis REGMODE_B="NOREG" */
           /* synthesis REGMODE_A="NOREG" */
           /* synthesis DATA_WIDTH_B="18" */
           /* synthesis DATA_WIDTH_A="18" */;

	 VHI scuba_vhi_inst (.Z(scuba_vhi));

	 VLO scuba_vlo_inst (.Z(scuba_vlo));

	 // synopsys translate_off
	 defparam sc_rom_monitor_0_1_0.INITVAL_3F = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_3E = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_3D = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_3C = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_3B = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_3A = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_39 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_38 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_37 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_36 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_35 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_34 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_33 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_32 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_31 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_30 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_2F = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_2E = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_2D = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_2C = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_2B = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_2A = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_29 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_28 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_27 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_26 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_25 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_24 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_23 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_22 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_21 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_20 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_1F = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_1E = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_1D = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_1C = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_1B = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_1A = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_19 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_18 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_17 = 320'h0000000000000000000000000000000000000000038FF034D2038FF034C2038FF0349A038FF03EFF ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_16 = 320'h00D00038FF034CA038FF03492038FF0348A038FF03482038FF0344A038FF03442038FF0343A038FF ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_15 = 320'h00D6300D5A00C5803EFF0136300D0302E0803EFF02E0803EFF038FF00D5A03EFF00D630105801363 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_14 = 320'h00D0302E0803EFF02E0803EFF038FF03EFF02E70038FF034DA0170801F100110801F100110801F10 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_13 = 320'h0110801F100110801F100110801F100110801F100110801F100110801F100110801F100110801F08 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_12 = 320'h02E0803EFF02E0803EFF038FF02E7802430038FF03EFF02E780110801F0803EFF030E800DE700AE7 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_11 = 320'h00AE400AE300AE300AE300AE300AE200D0000D0000D000342000D0000D0000D000341800D0001708 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_10 = 320'h01F100110801F100110801F100110801F100110801F100110801F0802E0803EFF0347000D0001708 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_0F = 320'h024700347000D00017080247002E08016E7016E4016E3016E3016E3016E3016E200DE7030E800DE7 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_0E = 320'h00AE703EFF010E003EFF010E003EFF010E003EFF010E0016E0016E700DE7030E800DE700AE700AE0 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_0D = 320'h00CE003EFF00CE003EFF00CE003EFF00CE003EFF016E700DE7030E8034700171002470030E801108 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_0C = 320'h01F0803470017100247000808030E80081003478011080081002478030F800AE700AE70340700AE7 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_0B = 320'h0344F00AE70343F00AE700AE700AE700AE600AE600AE600AE600AE500AE500AE500AE500AE400AE4 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_0A = 320'h00AE400AE400AE300AE300AE300AE300AE200AE200AE200AE200AE100AE100AE100AE100AE000AE0 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_09 = 320'h00AE0030F000AE700AE70340700AE70344F00AE70343F00AE700AE700AE700AE600AE600AE600AE6 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_08 = 320'h00AE500AE500AE500AE500AE400AE400AE400AE400AE300AE300AE300AE300AE200AE200AE200AE2 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_07 = 320'h00AE100AE100AE100AE100AE000AE000AE0030E800DEF02EE8016E8016E800AE8016E80000800008 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_06 = 320'h0000800008000080080800DE8016E802400016E802448016E802438016EF016EF016EF016EE016EE ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_05 = 320'h016EE016EE016ED016ED016ED016ED016EC016EC016EC016EC016EB016EB016EB016EB016EA016EA ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_04 = 320'h016EA016EA016E9016E9016E9016E9016E8016E8016E802600016E800DEF038FF00D0700DE702EE8 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_03 = 320'h00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_02 = 320'h00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_01 = 320'h00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600 ;
	 defparam sc_rom_monitor_0_1_0.INITVAL_00 = 320'h00D000380003E0002EE0016E703E0002EE80260000D0000D0000D0000D0000D0000D0003E0002600 ;
	 defparam sc_rom_monitor_0_1_0.CSDECODE_B =  3'b000 ;
	 defparam sc_rom_monitor_0_1_0.CSDECODE_A =  3'b000 ;
	 defparam sc_rom_monitor_0_1_0.WRITEMODE_B = "NORMAL" ;
	 defparam sc_rom_monitor_0_1_0.WRITEMODE_A = "NORMAL" ;
	 defparam sc_rom_monitor_0_1_0.GSR = "ENABLED" ;
	 defparam sc_rom_monitor_0_1_0.RESETMODE = "ASYNC" ;
	 defparam sc_rom_monitor_0_1_0.REGMODE_B = "NOREG" ;
	 defparam sc_rom_monitor_0_1_0.REGMODE_A = "NOREG" ;
	 defparam sc_rom_monitor_0_1_0.DATA_WIDTH_B = 18 ;
	 defparam sc_rom_monitor_0_1_0.DATA_WIDTH_A = 18 ;
	 // synopsys translate_on
	 DP16KA sc_rom_monitor_0_1_0 (.DIA0(DataInA[18]), .DIA1(DataInA[19]), 
				      .DIA2(DataInA[20]), .DIA3(DataInA[21]), .DIA4(DataInA[22]), .DIA5(DataInA[23]), 
				      .DIA6(DataInA[24]), .DIA7(DataInA[25]), .DIA8(DataInA[26]), .DIA9(DataInA[27]), 
				      .DIA10(DataInA[28]), .DIA11(DataInA[29]), .DIA12(DataInA[30]), .DIA13(DataInA[31]), 
				      .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), .DIA17(scuba_vlo), 
				      .ADA0(scuba_vhi), .ADA1(scuba_vhi), .ADA2(scuba_vlo), .ADA3(scuba_vlo), 
				      .ADA4(AddressA[0]), .ADA5(AddressA[1]), .ADA6(AddressA[2]), .ADA7(AddressA[3]), 
				      .ADA8(AddressA[4]), .ADA9(AddressA[5]), .ADA10(AddressA[6]), .ADA11(AddressA[7]), 
				      .ADA12(AddressA[8]), .ADA13(scuba_vlo), .CEA(ClockEnA), .CLKA(ClockA), 
				      .WEA(WrA), .CSA0(scuba_vlo), .CSA1(scuba_vlo), .CSA2(scuba_vlo), 
				      .RSTA(ResetA), .DIB0(DataInB[18]), .DIB1(DataInB[19]), .DIB2(DataInB[20]), 
				      .DIB3(DataInB[21]), .DIB4(DataInB[22]), .DIB5(DataInB[23]), .DIB6(DataInB[24]), 
				      .DIB7(DataInB[25]), .DIB8(DataInB[26]), .DIB9(DataInB[27]), .DIB10(DataInB[28]), 
				      .DIB11(DataInB[29]), .DIB12(DataInB[30]), .DIB13(DataInB[31]), .DIB14(scuba_vlo), 
				      .DIB15(scuba_vlo), .DIB16(scuba_vlo), .DIB17(scuba_vlo), .ADB0(scuba_vhi), 
				      .ADB1(scuba_vhi), .ADB2(scuba_vlo), .ADB3(scuba_vlo), .ADB4(AddressB[0]), 
				      .ADB5(AddressB[1]), .ADB6(AddressB[2]), .ADB7(AddressB[3]), .ADB8(AddressB[4]), 
				      .ADB9(AddressB[5]), .ADB10(AddressB[6]), .ADB11(AddressB[7]), .ADB12(AddressB[8]), 
				      .ADB13(scuba_vlo), .CEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB0(scuba_vlo), 
				      .CSB1(scuba_vlo), .CSB2(scuba_vlo), .RSTB(ResetB), .DOA0(QA[18]), 
				      .DOA1(QA[19]), .DOA2(QA[20]), .DOA3(QA[21]), .DOA4(QA[22]), .DOA5(QA[23]), 
				      .DOA6(QA[24]), .DOA7(QA[25]), .DOA8(QA[26]), .DOA9(QA[27]), .DOA10(QA[28]), 
				      .DOA11(QA[29]), .DOA12(QA[30]), .DOA13(QA[31]), .DOA14(), .DOA15(), 
				      .DOA16(), .DOA17(), .DOB0(QB[18]), .DOB1(QB[19]), .DOB2(QB[20]), 
				      .DOB3(QB[21]), .DOB4(QB[22]), .DOB5(QB[23]), .DOB6(QB[24]), .DOB7(QB[25]), 
				      .DOB8(QB[26]), .DOB9(QB[27]), .DOB10(QB[28]), .DOB11(QB[29]), .DOB12(QB[30]), 
				      .DOB13(QB[31]), .DOB14(), .DOB15(), .DOB16(), .DOB17())
           /* synthesis MEM_LPC_FILE="sc_rom_monitor.lpc" */
           /* synthesis MEM_INIT_FILE="rom.mem" */
           /* synthesis INITVAL_3F="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_3E="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_3D="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_3C="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_3B="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_3A="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_39="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_38="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_37="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_36="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_35="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_34="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_33="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_32="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_31="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_30="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2F="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2E="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2D="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2C="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2B="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_2A="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_29="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_28="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_27="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_26="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_25="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_24="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_23="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_22="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_21="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_20="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1F="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1E="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1D="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1C="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1B="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_1A="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_19="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_18="0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" */
           /* synthesis INITVAL_17="0x0000000000000000000000000000000000000000038FF034D2038FF034C2038FF0349A038FF03EFF" */
           /* synthesis INITVAL_16="0x00D00038FF034CA038FF03492038FF0348A038FF03482038FF0344A038FF03442038FF0343A038FF" */
           /* synthesis INITVAL_15="0x00D6300D5A00C5803EFF0136300D0302E0803EFF02E0803EFF038FF00D5A03EFF00D630105801363" */
           /* synthesis INITVAL_14="0x00D0302E0803EFF02E0803EFF038FF03EFF02E70038FF034DA0170801F100110801F100110801F10" */
           /* synthesis INITVAL_13="0x0110801F100110801F100110801F100110801F100110801F100110801F100110801F100110801F08" */
           /* synthesis INITVAL_12="0x02E0803EFF02E0803EFF038FF02E7802430038FF03EFF02E780110801F0803EFF030E800DE700AE7" */
           /* synthesis INITVAL_11="0x00AE400AE300AE300AE300AE300AE200D0000D0000D000342000D0000D0000D000341800D0001708" */
           /* synthesis INITVAL_10="0x01F100110801F100110801F100110801F100110801F100110801F0802E0803EFF0347000D0001708" */
           /* synthesis INITVAL_0F="0x024700347000D00017080247002E08016E7016E4016E3016E3016E3016E3016E200DE7030E800DE7" */
           /* synthesis INITVAL_0E="0x00AE703EFF010E003EFF010E003EFF010E003EFF010E0016E0016E700DE7030E800DE700AE700AE0" */
           /* synthesis INITVAL_0D="0x00CE003EFF00CE003EFF00CE003EFF00CE003EFF016E700DE7030E8034700171002470030E801108" */
           /* synthesis INITVAL_0C="0x01F0803470017100247000808030E80081003478011080081002478030F800AE700AE70340700AE7" */
           /* synthesis INITVAL_0B="0x0344F00AE70343F00AE700AE700AE700AE600AE600AE600AE600AE500AE500AE500AE500AE400AE4" */
           /* synthesis INITVAL_0A="0x00AE400AE400AE300AE300AE300AE300AE200AE200AE200AE200AE100AE100AE100AE100AE000AE0" */
           /* synthesis INITVAL_09="0x00AE0030F000AE700AE70340700AE70344F00AE70343F00AE700AE700AE700AE600AE600AE600AE6" */
           /* synthesis INITVAL_08="0x00AE500AE500AE500AE500AE400AE400AE400AE400AE300AE300AE300AE300AE200AE200AE200AE2" */
           /* synthesis INITVAL_07="0x00AE100AE100AE100AE100AE000AE000AE0030E800DEF02EE8016E8016E800AE8016E80000800008" */
           /* synthesis INITVAL_06="0x0000800008000080080800DE8016E802400016E802448016E802438016EF016EF016EF016EE016EE" */
           /* synthesis INITVAL_05="0x016EE016EE016ED016ED016ED016ED016EC016EC016EC016EC016EB016EB016EB016EB016EA016EA" */
           /* synthesis INITVAL_04="0x016EA016EA016E9016E9016E9016E9016E8016E8016E802600016E800DEF038FF00D0700DE702EE8" */
           /* synthesis INITVAL_03="0x00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600" */
           /* synthesis INITVAL_02="0x00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600" */
           /* synthesis INITVAL_01="0x00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600" */
           /* synthesis INITVAL_00="0x00D000380003E0002EE0016E703E0002EE80260000D0000D0000D0000D0000D0000D0003E0002600" */
           /* synthesis CSDECODE_B="0b000" */
           /* synthesis CSDECODE_A="0b000" */
           /* synthesis WRITEMODE_B="NORMAL" */
           /* synthesis WRITEMODE_A="NORMAL" */
           /* synthesis GSR="ENABLED" */
           /* synthesis RESETMODE="ASYNC" */
           /* synthesis REGMODE_B="NOREG" */
           /* synthesis REGMODE_A="NOREG" */
           /* synthesis DATA_WIDTH_B="18" */
           /* synthesis DATA_WIDTH_A="18" */;



	 // exemplar begin
	 // exemplar attribute sc_rom_monitor_0_0_1 MEM_LPC_FILE sc_rom_monitor.lpc
	 // exemplar attribute sc_rom_monitor_0_0_1 MEM_INIT_FILE rom.mem
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_3F 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_3E 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_3D 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_3C 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_3B 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_3A 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_39 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_38 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_37 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_36 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_35 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_34 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_33 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_32 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_31 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_30 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_2F 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_2E 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_2D 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_2C 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_2B 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_2A 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_29 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_28 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_27 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_26 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_25 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_24 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_23 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_22 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_21 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_20 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_1F 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_1E 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_1D 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_1C 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_1B 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_1A 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_19 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_18 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_17 0x00000000000000000000000000000000000000003FF8C300003FF8E300003FF90300003FF923FF5B
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_16 0x1004F3FF95300003FF97300003FF99300003FF9B300003FF9D300003FF9F300003FFA1300003FFFB
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_15 0x0000130001100003FF691001400000068003FF7E058003FF803FFFB300013FF7800001100001FFB3
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_14 0x00000068003FF89058003FF8B3FFB93FF9B008003FFBC300000FFBE1001B000331001A0002C10019
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_13 0x00035100180003510013000301001200030100110003010010000301000900030100080003010007
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_12 0x010003FF97058003FFAA3FFFC00800078003FFDB3FFBD0080000004100063FFA2000000001C10004
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_11 0x000083000C2001010014000183001C0000000000000001000000000000000000010000100010FFF3
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_10 0x10063000481004D0003F1006D0003E1007200024100570001D10077010003FFC210000100540FFFF
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_0F 0x0080010000100540FFFF008000700010004000083000C2001010014000183001C0FFE40000000008
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_0E 0x100043FFDD100083FFDF100093FFE11000A3FFE31000B10008100040FFF8000000000C1000410008
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_0D 0x100083FFE7100093FFE91000A3FFEB1000B3FFED100040FFF400000200000FFFF010000000000002
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_0C 0x10054100000FFFF01000100FF00000100FF000000FFFE10100010000000000070300803000030090
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_0B 0x300003008C300003008820078100743006C2006810064000603005C2005810054000503004C20048
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_0A 0x10044000403003C2003810034000303002C2002810024000203001C2001810014000103000C20008
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_09 0x100040000000070200802000020090200002008C20000200883007C100743006C200681006400060
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_08 0x3005C2005810054000503004C2004810044000403003C2003810034000303002C200281002400020
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_07 0x3001C2001810014000103000C2000810004000001F9940E000000001007410000100841000110001
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_06 0x100011000110001100FF1F99410090008001008C0080010088008003007C20078000703006C20068
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_05 0x10064000603005C2005810054000503004C2004810044000403003C2003810034000303002C20028
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_04 0x10024000203001C2001810014000103000C200081000400000000001066C3FFC530000007F40E000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_03 0x000000003B000B500800200800000A00000000000000000043000BD0080020080000120000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_02 0x000000004B000C500800200800001A00000000000000000053000CD0080020080000220000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_01 0x0000000081000D500800300800002A00000000000000000063000DD0080020080000320000000000
	 // exemplar attribute sc_rom_monitor_0_0_1 INITVAL_00 0x0000000091000E500800300800003A00000000000000000000000000000000000000000003F00000
	 // exemplar attribute sc_rom_monitor_0_0_1 CSDECODE_B 0b000
	 // exemplar attribute sc_rom_monitor_0_0_1 CSDECODE_A 0b000
	 // exemplar attribute sc_rom_monitor_0_0_1 WRITEMODE_B NORMAL
	 // exemplar attribute sc_rom_monitor_0_0_1 WRITEMODE_A NORMAL
	 // exemplar attribute sc_rom_monitor_0_0_1 GSR ENABLED
	 // exemplar attribute sc_rom_monitor_0_0_1 RESETMODE ASYNC
	 // exemplar attribute sc_rom_monitor_0_0_1 REGMODE_B NOREG
	 // exemplar attribute sc_rom_monitor_0_0_1 REGMODE_A NOREG
	 // exemplar attribute sc_rom_monitor_0_0_1 DATA_WIDTH_B 18
	 // exemplar attribute sc_rom_monitor_0_0_1 DATA_WIDTH_A 18
	 // exemplar attribute sc_rom_monitor_0_1_0 MEM_LPC_FILE sc_rom_monitor.lpc
	 // exemplar attribute sc_rom_monitor_0_1_0 MEM_INIT_FILE rom.mem
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_3F 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_3E 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_3D 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_3C 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_3B 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_3A 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_39 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_38 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_37 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_36 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_35 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_34 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_33 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_32 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_31 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_30 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_2F 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_2E 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_2D 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_2C 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_2B 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_2A 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_29 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_28 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_27 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_26 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_25 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_24 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_23 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_22 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_21 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_20 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_1F 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_1E 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_1D 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_1C 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_1B 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_1A 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_19 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_18 0x00000000000000000000000000000000000000000000000000000000000000000000000000000000
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_17 0x0000000000000000000000000000000000000000038FF034D2038FF034C2038FF0349A038FF03EFF
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_16 0x00D00038FF034CA038FF03492038FF0348A038FF03482038FF0344A038FF03442038FF0343A038FF
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_15 0x00D6300D5A00C5803EFF0136300D0302E0803EFF02E0803EFF038FF00D5A03EFF00D630105801363
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_14 0x00D0302E0803EFF02E0803EFF038FF03EFF02E70038FF034DA0170801F100110801F100110801F10
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_13 0x0110801F100110801F100110801F100110801F100110801F100110801F100110801F100110801F08
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_12 0x02E0803EFF02E0803EFF038FF02E7802430038FF03EFF02E780110801F0803EFF030E800DE700AE7
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_11 0x00AE400AE300AE300AE300AE300AE200D0000D0000D000342000D0000D0000D000341800D0001708
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_10 0x01F100110801F100110801F100110801F100110801F100110801F0802E0803EFF0347000D0001708
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_0F 0x024700347000D00017080247002E08016E7016E4016E3016E3016E3016E3016E200DE7030E800DE7
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_0E 0x00AE703EFF010E003EFF010E003EFF010E003EFF010E0016E0016E700DE7030E800DE700AE700AE0
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_0D 0x00CE003EFF00CE003EFF00CE003EFF00CE003EFF016E700DE7030E8034700171002470030E801108
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_0C 0x01F0803470017100247000808030E80081003478011080081002478030F800AE700AE70340700AE7
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_0B 0x0344F00AE70343F00AE700AE700AE700AE600AE600AE600AE600AE500AE500AE500AE500AE400AE4
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_0A 0x00AE400AE400AE300AE300AE300AE300AE200AE200AE200AE200AE100AE100AE100AE100AE000AE0
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_09 0x00AE0030F000AE700AE70340700AE70344F00AE70343F00AE700AE700AE700AE600AE600AE600AE6
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_08 0x00AE500AE500AE500AE500AE400AE400AE400AE400AE300AE300AE300AE300AE200AE200AE200AE2
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_07 0x00AE100AE100AE100AE100AE000AE000AE0030E800DEF02EE8016E8016E800AE8016E80000800008
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_06 0x0000800008000080080800DE8016E802400016E802448016E802438016EF016EF016EF016EE016EE
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_05 0x016EE016EE016ED016ED016ED016ED016EC016EC016EC016EC016EB016EB016EB016EB016EA016EA
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_04 0x016EA016EA016E9016E9016E9016E9016E8016E8016E802600016E800DEF038FF00D0700DE702EE8
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_03 0x00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_02 0x00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_01 0x00D000380003E0002EE0016E703E0002EE80260000D000380003E0002EE0016E703E0002EE802600
	 // exemplar attribute sc_rom_monitor_0_1_0 INITVAL_00 0x00D000380003E0002EE0016E703E0002EE80260000D0000D0000D0000D0000D0000D0003E0002600
	 // exemplar attribute sc_rom_monitor_0_1_0 CSDECODE_B 0b000
	 // exemplar attribute sc_rom_monitor_0_1_0 CSDECODE_A 0b000
	 // exemplar attribute sc_rom_monitor_0_1_0 WRITEMODE_B NORMAL
	 // exemplar attribute sc_rom_monitor_0_1_0 WRITEMODE_A NORMAL
	 // exemplar attribute sc_rom_monitor_0_1_0 GSR ENABLED
	 // exemplar attribute sc_rom_monitor_0_1_0 RESETMODE ASYNC
	 // exemplar attribute sc_rom_monitor_0_1_0 REGMODE_B NOREG
	 // exemplar attribute sc_rom_monitor_0_1_0 REGMODE_A NOREG
	 // exemplar attribute sc_rom_monitor_0_1_0 DATA_WIDTH_B 18
	 // exemplar attribute sc_rom_monitor_0_1_0 DATA_WIDTH_A 18
	 // exemplar end
      end
   endgenerate
   
endmodule
